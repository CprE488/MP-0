XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x<��!�	oЗ�Q����܉�I$
��ĥ���Ϡ�wŢ�d*�@��礰]��
LG�:|9)��G�,K�K���g�=�n��Hw9�˛� ��~%� 1�v<�Ǒ�����3f<��vߒ _�Ե�-M����ɢ�����,`��c���m%!X��������U�G�D�Ԭ��TK�Yb�+'�mj������t�Y��ϝ�;�&Y)3Z��ة86,��F�4�k [���]����Lw�U�5#P7��ki֤mH�T�F����{!jǅ����Zi�r ���T)<�+��V��8���+W|�5�+ň�.�����4��V�d �k������r*��?����4��%�Y�?�2�5��S|�mgj�\pÒ/��2r;/��:
���"; .x��N���C2q����Ha�oY�9�wF��6u��h{�"�i)ڴ.��pyGUh�����h�������O��)���}pR"�ܓ��)X��{ɚ2
�����[����i��������<w~�BҘ~q>�~Z��p �<9/M���l�׍���اF "xuC����,�Q7��,~�Ϩ�����h<�F$��a1�]vo��Կ��{	p<W�J4m�!j�dr�����)V�o`�����5��q��UmC�*�����M[a�M�4H��j>k�� hwT�C�3w�3�o�T�%<[�����	m��`~��
\�uCD�զZ��s�Udv�?&}�o�.1'M )#T�����Z>f�
�"����e�=~��i�:��XlxVHYEB    95d3    18d0������
�W!��s�eof�N�cL��#�܆J��
ֈ�@������8�J�	*�	�m���ٹ2Jb�	8�BbY!]'�gwhf�I�$w��$��o,����:�읫��{2`�PK��? ,dXi�d��t>��`v��h!k�թ�,2gr�DA�s�Ct�~Kg7�JZ�a9���>/�������R��G�ӂ���E�.�JѽϮ�	I^��^��5��Z>�z~�/\��`۷�d�)ֹ3h����?|�j^�7��������8O��V���P�D.��K�Δ��A��T u�ֻ��`3A�g������"Րm�R�v�R�XTJd�<8��	.9��L��8����b���o�x����LJ��_�
O�uV�-e /N=i��ո�7�3�Wה\�m�'��}p	+���t�mшP.��3�G�u���1�hL����o:�,f��[�*� ��������~��%;������ֻx���Q1��!��+�m�ߤ���R����Z��S�wo�6�팔�Wh8�k6~�nDTm�G�S����y݊v/6	����|�b���"��!�A�EZ�'������u�$�n@d_$����CV[��i�m%O�+��2��kQ����u��q7>�J�
���cp��������CĽS'��.l�.}��SjspĤ`�y�����0ǣ�P��v�^=\��7��۔G>d���C��^21�+Im$䅧�`ó*�u�D,��ǔ�}���B��t�����)3�L�rP"/@'���i@�Q.�Ul���8�MHE
��{�7R	z���@{g�Χ�����pԊG����]]��9g� f�f��C�s�H ��]����)�Z�1���S��:y�XX�Նs�\����ے]33`��o�ou���V+��7T��Ô\*������3����Cv��!j�zфfm�τz�t�A��]X�7搯dN����R�߼"h�(�;S�;���E�Z����}z��;�����!,L�����T�L%D}��&��d�x����^�)+:�/�7�����#X�a������.Q���ԗ�F#�rS����A��xVձs���^����XC�SU]E/������4/�@(.����*��C����Ɔ�F��Q�X���\�������/T�����
m�:TN���>]W��-�&�z�]Ӷ� EM]B��g-��	�jF����o���`��R���-v�� -����b���Z���S@PV�%�߇����C�h[� ��s�潹񡻈H]�<�)1�n^/ƴ���c�r���U�-<z�� 	�7�/H`{П�iI6�F�^O�ep�����d�@�I"�
�b0j��Ҟ#Jv���^t�b���Y���ȣog0*
�m�_0�e�C�/A:�7&���/M�z!�A���O!I�> #1���9����TU3����R�C�	��c�� a,�5	z����7������&����0�z�Wp�,�v �B�U�ʅ�㘟�DF�g�m�����3��?����Է���K�����Y���쀝;R�B�����S୨�<G[~��R�����p�BI�ΐm/g�$���_�tLe��9=�=d���U��4�1��O�����.U�3�9�^�� -�>��A�o�FU�Mǵ� ��p�D�]�c���YL�͔�%���Js*wn$ :�|�O���` �aێ߉- �*�j���e����5�IR|����kp\)�F�6�&�R-&~Kʡ��A��Z��pE�`;�_G��ވ�J ��zz�����B��X|Ű^6л>7Qd�vzB��g������;'%%��1rӄ�"�C�W�lI�S�$ecQ��y�&]��b�$�a:g A�/g�;>�sg
�������H��-yQ^�d�p�69mI�RKZ����SM���lY��	����E$������9b�R�����g�<ښ)8$�1��W���*n���y�V8[���q)�$�A��,�X�t�]�'k,MO�����XTQh�'�rC�e��% &d`H�s���s�٠�;��Tπ��|�N�asxE����]�۝��D�v���z���tBD�Y��O�f�Җʃ�\!"��~����pd�dv/���%�u<�B��n��Ͱk^/�ɪOS�ᇸV�.4̼���E����s�k�*ޛ���G^�0D죜r����v\+��z�1:�A�f)�( ��Nv(쩯�'�{z��8;���A���,/F"eЁ��F
'q���ơ �p�ö)OJ��y/C���r��iaD��$�,[�_*^�lI1X(S.b�[��@O��w�A���4��Dl�owI*��ў���%�ޣ*�z���r��S��Z:Mk>�U9�R�Ў���1�ӛ&�^���:A)�F1{:n��/�Ý��Z<Tw	��(�#�����?I�cne���_�X&JMK�ݠ�2mT���p��i\�=`Jٖ��F�Ml����N��"쀟�-.A�.�w�&1�K#5���1�=�*��ϒ���Nz&J2қe����P4u7O�9i�I�F�()'j�V(m�C����ÖO�"����-��8[�9"�@cZ�r�O�p!k�쬊f4ƞ��c#�緌��C=/ib^&DYAkR7��H6I�/�֤��6Q���BbP��������LH�Oq�bMz��y���O/�hv�/��B�qg�d��X���ޘԜ���S�]��b��\^Ļ<�8ߙ%�0;)���e������Y��'�?��uD��.��JRx
|2��)�6$Ł �Zʛ�cD��z�@�+7*x�Y�%�'D�<���wݨz�`�}��T���K(�/���b����~RT����'�z�}MSmP��nmgAӏ�6�������#7L���9� >F`�#*��*��<����O�$�T5n@TWM)A��!0��,���O�,�����+U��#��]H8�+�0o��bPY;�2~"�x�{��牥�n|�"u�Ô��p��O���H7w�q�]��/q��o+u��۳P�-�C���]N�c?��.��PJ��ZJ��8cH�MցQ�RM�]2�#{��If�����Մ.�ϜO�a���|K�[�[���*/AQ;�Uã�����ˁ�z �W=F ���HVN�_�5� fk�ƙ�j3H%�S�bT*���^מ������b���o��~@<C�z�N��h�bi;�Q��t;�.*�"
��8!������U�{��t�$�Cz�7���)���� �q�������V�����q|f�uo%�@����z����R�=����m�{�ܱ���t��2��������v@Z٬��=�W�E���/3��LcU5{��
�"o�[I�dY>a��+]����!�C�9�
#�㘪;=�e	.ǌ#�����E'���H�U�#@������/$��UwA��Ap��b�R_��B�C�7����'GX3��0��v�%�|U�֋ʒE�r�Y%x�fU�P�J�qR�ko��R���,�����Z�L��ɦ2��9��h\H�����j(3�Lh���ЉC��������%�7�EV�!��՜����x�3ka�O�e�Y���#8�V6�"	T[h�;C��~7�ZE5���`#�JYSJ�u���oAgj��ˊw�l�8��j,3��������٘pܭ^�?�g�] ��	�"~H��=i־�Ȱ7�R!���%kfa��dU(3�V:\�,�xq�v���Ǉ�����y$W��o[X�Eʝk�D�����4Ti)p֓M����vs.9^-�-_׃��s�+ʀ���2e�ܳ��.�c�=�\N�f��ǟ���X@��������EK����Ku�76I��� ���"�i��O4�>��	�m�����욤��1�"����&ݭ"<=��^���m�dјGIJ����̬�nb�|�	�V�1���N�຺$�m'�0NJ#�"='C���⟺kq���R'�ԧ;���y^pA%Lk"�lC�P�Orx��ހ���چv��'���8�.D��Ʈ���wƓ�!��9>)��}�;���F�eA*���_!i�t,���6r��~Ƽg���._��m����d
��`�s��D�E���[i��{D�!/)L�V�[.��@�s$@ӦہMF-�0�6���p���:x��f(=�,�	����S��]�W�k�ⳏ��]a��2���e��`%"s���q-��TH �[�ol8�nZo5�Du�)�3��%k���a����ݞ~���2�%��ݮ�>��; +�� �0��	�.�?���$0��I��p��0`�⽩�|�����-�O��s�p���̵@��>׀�4�\b&p���#�q��H$�$"����g�����c$�2%N�`9��Wئ>���k�h�b�M6��ӥ�e�#K����()�"��Nߑ7��?o��Q����=�O��ta_����0�j���o~�r�,�����KF�\�y�p� �$;����0t�_y�3z+V�a�d��1P�u�ë5��gJ�s��G��k=���9����t�J�H����3suː��D��_�e�@UU˨���/QC��,	�^���:ʜ����=�I���h�z�!N�����Xs�'T6L[������Pi�cl��l�srh��_��S�T0��E�80��y 0��N�5k�=�W���t�����\�B��V�Y���h��f^E�.�V��C
Hv���j�r�������n��9�3�:sݙ��;�n���6�:��(��9-*C��~�ڽ��/���2n�B�1������Q�����S:���h�ܦw�j"��� 5��A��G�(qL<�H0�02����t]���;O�����(3�Y�C�}�\T_8 w�~���m�;�ʔ�|BB8�pw
�ZO��+(k��B���J��\�P����A�-e{�L��u�����@��眚���Q�/}^����Np[�X Aܬ�  x��ʪX�t�������ߗ's�LUү������93Siٔ�u���9غX��6I}"��A��s�g����һi� l�?eб�7��l8g��>o/��N���N�,%��~�f8v7tm 1��Ӹ���CoܯV��ΗjÙų-�g�=���V����L���ᜁ�r-@�`�4\=n=�l�)�Y���O\�~ͭl��0*?�D̍_�r�NFMIm����&!r?��+��'%I�r>äR�-2&U�i ��<G*�T ^S�o%hA��Sz� '���=ݞs$�ݿq,�a�dW�0�%0}
�+�yR��؟��� ��� ��I�1~$$��^�gwG�X�k���r�5���KcZ�{
�+W���0|/��j5(:H������m�صb����a�-�E�������Ĉ���rޛ���eÇ�Z�A�ޓv4W<8�U�Ra U�F�s'��հ�t�~�}�)h=�Zmaʱ)�w^
)�������.#���tIJ>��8����L�����%TwO�<R0ВΘK�G�)v���]�	�i��^�U�[����18�Q^< �n���+��Z�����Ȭ�p2!&��Gn�_���r�'#��Δ�W�OQ��y���k�Z�F ��޸L@_\Q@K�����346�y�;lr�#>Y������	�VK��Ƭ�Y�x��yW��FHD#iRn��]9Ƥc����G|P�C��gP���뤓�Fb��!�'��D:Ic�^ӆ�bQD,[�Yq�alJ�-C���ӆХ��EY�G� Wi�����!���p�v�/�x�]��wovˇ�R�HhiҌb֓*�^���f���=���r�U&*@�xA��%o6�|v@��vc�H���4���S���S�ؼ�E��j"�G�.>�7K�T��`E���W.�Fr{9jd�3n�OKOD���|k�r�p�V�a(�(-�����''�myY]Gx�$��RW�n�]a��<�<��U�|��:�M�?���itN�9����L+8W�zg5��!��+�p������00�.�cbA�<oJ�+���=�%��'�ϴ��>壋�xX���)���B����
���_'>���p�<p�쒼S��
Ǭa�S< ���qvo���)�tI��dQ'!:б��#�����QS��ݙBl��O;��Q�^J�C�ɭ�˸ڻ��EC3 2�