XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]�+�Ԏ���~+�q�!����ޙ�  V�0|���eb�D�[�V�LX��2avx��' �/y���¢^�s�XW/�*cU@&�����,�]��i��>�Ж�Î�&iY�*Jn�b��{�U��|���+���C�T�a��F�N�lj�`�nL�1i;��r���>~3Iݗ����F��cU*��������SN-��<%�
��,���lMn�m��E�R9լs�������9����B|$���`g�!_����DL�Ҝ<:�e�^�d?,d���ף�!V(�h���տ7�-�%�Ā2Us�TX�n���sVQZ�ـ"��HIP�*�oz��Wlmw���O��6�闤��&���� ��%����5��L� ���ر�B������IC�ϋ��+]�����L3:�k�zG����d������|\^62B	��+:_����%�&��Z���kzX��4Q�BH��2:~�n�u3���e_���:�������Y�;4e�}�x����|2�f�u���+������a�m�{���To
����	*�;��W�X(���w���hS�2X��*�%G�ʮ���ϠܼQ�y�S�؁ШJ�K+u��J��aR����������vn�UJ���x2;�]q2�b^z���yYgߴ�/�,�Y;T�2�Xa��B��M�˙���Տ���Z~��hb��l� �s��4��Zx��(E;m��(�ꯨ���!-O���XlxVHYEB    dd8f    2160Vى}�ЛslYxE7�Fb`M.�o��,e��q�5AC���0qk���(��� �):Ƹ�Et��@)C��mI>m��Z���r���W�G�7&����f�Ʀ�d1i�T~����޾�JK����
��EH{�u�8���@���	R�:���L����zb9ڋ$9CI��E�1p!֨�%LN��K�h����ˡQ3*��p }��ES�/�0s������F�f�i���Ճ��1ӇC륓j��#kJo$�]/�u���Tb�	Y��:@�7����ܳ���OXa��]��j����d�w)%��v�`퓂�����c3�R���:��Q�D�0^.��j�?F���xdupk�|����3��RMy��O�i���,x��s��|����r��
�W4Y��V���*���זSd��ɊM�Ԃ`�G�h���c�$��^�����9j&�6zy��P-�3"�R�:w$���$o;P�p������$���V�����Z5���^�������b�8\M�I�׃M�����֤8\CTGrv+����c�>i�-1���B�^�8p rO1�.�'�t ��W�n���س���,�aOTg�ڬ�e���F�y5 ���BdL�oې=�{�ԙ�  �N��2�UZP@�d'�g���jЁ�4�y�~LXLw��'�<>:G$�N)��xbn8��,,���n�?-�f�7���l%����#/�?�}��H.-�w�Fg%�o�hM��(a^��M�9y�u�K(�&x68�h\�.]',$U���)qB�&��s���P���P��T5���Z����. 5y\e�������}=�.�!�Z]w,V��jv+��Q�&�@@�?q��H���G��G�y]& پxH^e�c�������Z�3����!��p�c�A�ux�&�\���kU�팿p��	����j�^�<���/7sm�pΔ,H7�ީv�[HkLV=F�J����}�
���?��(�km�G�-��)p�&VҩQ�q�\��T�3t���\��|ب���� ����� �B�߁�T�2�YsP�0���*����7�'��qW�o��JeО�"b�dܗnt.�*���sy��9|�	$a���P&�I�э�>��S�@X�&2[�*=�TEd�Ec��X}c�;I&<UO���m;�.(K4_(5�0/,8B�H<.{��O���_p!>�I
K���h@xM�|��=�e����&��|�A;|&������/���v�xގ�N�C�,�R�K���veZ�����nN7{4��XGJ��2[�n$:& ���^䀊����3R�7����m��{��$O�o 4���ҿD���]�r��ޙ)̄��kg����;�F)����1�P����w�q:Z���q�J�:�!��G�^d��o����v�V�2�.� =�\Q\�4������`�xԻ��h��מ���S��
@��m�rQ��c�������K�m#2�l��J�H{��U��4R�^hK���N�eJiv�l ڧ��*+/��T�D�`���&j}���1� M���Z�<_�@lZ2\"�:��/����y'F�>BҜބ�F�]��@S�-�� 8�dQ���w�́z�~�yk	�h���G�
fi,�e\W^��A��g�����7��90*=629��8%j��i�^�E��m�!��)z.`G��o �ZK�aw�7ݹo?*�mtb����m~�����z1j�aD~=��iҭyH͑w��i֛V0���fn��}���*w�&�D�ap˼�p�\���$���x�Sr]�r3A$5��J#x��f��_���V1�5%s��F{�M��* 3W���E���u�d҅� ����Z���"�J ,�&#~Nw��j�+v�Z�9�Ƞ�`�w�{h<�^\���ZR�$'k�P ��$2���h���Wn[��&r�G��Hՙmp�[\�ڇ��O�B^�	m��o��lНBǘ�Hs�}�ϘN��S����kO���i�S�+H:՘F�Ͳ9��E���O����b2��L�_(��Р�y�{qFN0�.�JV�#-*�9uD0Ӿ�W������&R�M'�C��=A>�a�s�8D��X2�fV:�#�����oXz[���4~@�4��.�9��j"��F�K�e*�f�N_볃�����S���'q9��2��6\�PԠ��9���pv��\��	��!��UnD������?i1[`���w�ժB�Q��"B:���hS�[�ms�n�O��T�U9�!Ҁ��{��qa�w�z�8��%�0��¢�nY �}�?��X¹�hT����>�V���@`6 "�b�:��;�jxN}Y�E���q?Rш*�:�y1����p����κ=�ڗ4/K�|��VWtGe�x���wt-%�P����#�QD&G=%�fBw��p�H�yP�G�c)��:��:�n�!v���K�#�4#��f��� �����7���[s��@�K�����޴��*�̨���0_o�b���F��sjN����^@J��Kvc�1Nk�oQ>��~0��̰*�2�<}���"���Q�Y���Ӈt[dV�gF������f�-W�&�z-�F�XCtP9���&���67ަ!Rkz�js_�Ҫ�m��ۤ(.�*�F?�ʳ�{&��Nz�2�X,T��Q����26�#fTǇ�_�)D����TZ	#F6 �>�À�]�A#�Ln��RZ�@Y �Sm
�]�����`��El�X}�l��Ԛ2f�����b��<N���2^X�ŭ�O�~o�������զ�(O{aC�;�p.��Ἠ[8j���wv�u�Cf
�z����v��% R%�7��:���Wy
�U/.��0xE���14~��ʤC�y��5ok��r�]͝GɃ���F\ؼ�CGA���d���}� ��{o&�yO� �RI��2X�CO���� ��C���.�?�����j�v!���E�4�`��f��U�E~��9R�Y�S����YG6qG��R`xu~%����u���]�ë�1p�eT����-�t� ��]J�3y����M�=[-�'�]��[��#�N�f��"G���6��C&��OlGE�CdDJ������N�E\�����Y����@3�������^�SS�5s��5���F�*���X
l���GX]C�����'
� ���9pe�<�{v��� ��G�Ǿ>b>���P]�����7��E�CԺ�f�*D�Ro�7V����G��x�#xzs��F�&�ee����p��=T�F	ȁ>��2 �8�"��7U��3����м�z�F$󔃓�v�p��2�Ő�aDN"u8G�G��՟���R�naZ-j|��q�R)��"k�+D���V����=)�!�L`�5I�}�Jg��G��=�,�2W�r%�n��<��>�I����.�6m`��0�+T��JΪ��4�GOx�&}�@���AX���y�qǪ[yP�+g���>���� @�5�"$ԛ�f'
�
QP����|�z��b�'��$h��!/�ؓ���IM�Eh}�� �96���o�����5A����x�� �W�?*�uf{�Bp�1��	���B�;,H��jz� ��_���rښ�OSS}>��3�j����A&�d����W�I��`Y��|����:*_�33���3h�Ӹ�C�����a0*�~���b_���uU��V�����
��:߾͛J�`�z	D�.{�ǘ���� ��o�=�> ڍf	���3?�ݬ{R�i������cv�0���j#����d����h�a��d�n&��1�!�8�rv���~� ��B�|_�j���e�4�1��w�f��>�ښ���[�ڴnd�5م鞊��j~	.�E(e�lQpS��[ޫUr	���}��󢿱���.��yyyh��O�깣.ZӢ�Z��>&:lĕ�T������j�����l@n*�O�8�{��=��3�@^s�x����u�D�1�d�_�%������ U̩[޲�;�L�p�n1�&+�;�,.U�v�l�Q��AB�� ��a�%wS����3��%ob@���/��l���9�&��1D��]QL� ���v��׌zme���9!}j2?��B���61���,����q�;�Z��^�I��J���[�v��4�H���&-y�[UW�k�R9�"�;* 1�FӈW���ʘ�Grp��@$�-x���R��������A��?��I4Q�/�t�̟��5��ߗ�&�ɩ��I�=��.Q�f�$F�&��SY2�0�f�oW�����U��:�[��aDȇ	7b���ɂB�u�o�B����oC<�.�te~���.[�����\����6q�ϐ^�ѷ���\<L�5�P�
*���>7jbTG� $W3�:kUemkO�G�7U.]��"2=���&�ԕ�\�r�k7;��~���S�i��t�]�uTϷ
�HtB6y{/e�(td�V_��u�Q�$0t��<�	{��8��'P�;`)��L�+
J�������M���^]+���2,��<e� �+8��2A�j�5��v��) +�)n���ݪ�ͳ9�C�ۊ�w���1��t�KP���(��kfd1�ɺn��i-e)�=z�����D<������9܈������\>�b�_�D7�(�$;&�T�0���ӹ^��(������gXR��x����qA��B廅����R]�W	a���<OA�b�`>�8��d����P��`��*I��!��вJ؄�OMj}�[�)���\���]�ڻ�(<o�eS�6˘�"�D,�_��A붼Q�ES�̸W����&y��џ��ޱ�@���cKM�?Y��}O� �ϣ��ս�:���=�+��	�{�PB��EK�˚��HF�m��<�_e�os�E*�h�<1~������`�.P硅%?��b�!�z-ǚ(�r2'�R�!��
�
��M�E�_B�r�D߯��x��������z��D�Z5�zv(��Y����f�>�U��Tk����zr�[�<�:}Aa��U��(�J7���۵3�P@���u��&j3���[����SkJ� ��It@�tÒ���I���������{��L��$
��Y�ȿZf�|�]��0���<L�|p��k2�<t�N���u{e��m;�SO/�
 �Y�a��	⃘ `φFU�7�T,���v��U.p��׏�J�;LW)D��:�����7�;�����࿜>�G��w����(�ҥ�`3p<y}׍�ܩEFW�����+�"���3<��sQ���5<�w(7�j�l{���6F�C3�ZZ�݇�[ zV��H1�5b��P~���ប��B� uc�I~R@�����N.'t>�]�?GN����tO�;�A{�s3R]�O�S���eL~�5�� �
�z�5O�W��J�'\�Q6�D� Xd��I�E8q{{�e���BT-�΃M4�G�� ����~��Y�W���4���:ƭ�ЕF1<5�9�S���':ӏ9�oЯ!\�e;��/lL�䂭���c�d����F@��#0ȯI.%�A���=�f I�żFŤ*��Ԃ�z�24.Jj�ق�h
��Y*��X5��RdG�A����۲���[Ls� 
`7{XT�V�3�X�\�B���_=���N��,7��s6�{�ȣ��{�z ˅�H��G������5�I؎�1���$�j�E�F�D�|"��O�T�Ŗۏ[�Lũ���N�6�V>��%�{��`N(�S�����=3.PU�|��'���F+o���)�H�]I�(]�M�^`-��:���V|b|Y���8���R4�P �_paL�n����u�F'�׸�A����d"��7oӱst�4���J{Y	g��&v��P�V�K�T���4�T����%�Bk�es�0�7)p��y	��D���Kf�0��NZ��.K�6�ڔu�8 k�°e�:��ƞ
3���7u3�(�*&!��;���#��X%�y�m~�����m���Ժ���̓�C��d���_�톱4Z�t��r�?��$`��jTnb`�����I7'�Ċ�	4��)Ljg��r��� &�Cu.6��4��)t]&W��b��f���&��Ү��� &3]))�QS�C!���u��_�U��B�d����K��Y�ߝ��d��ϥh��%���wU �JcƄ�yc�=�j������7È���s$��X�����	�qh���7;�R���`FH�B-I��y5���Lr^�o��ϵ�TgT����Lr�/$s�ˏ���{?�glH��!��0��僑� `_���~9{t�>wJjv���D��Ǥ"��${���C]:�o_r?#ﰑ�[Iz����R�@��s+��H�:C���~g7���a�	�2O������d	�u�X����Κ>�5l碤!�o�q�\�����������e�`$��B���s3�J;�"o�u�'`F��D�����ק��ɗ�׬�)L�I�[~���8��i���uϾ] Ɣ�W���ȟЈl1��{V��**��7���F��D�i������87(1�Ϝ�K���5o�2����<0LU��Z�j��?|H꺌����kh�4��i��Z�r�Qe�oX��b���"srY9����܈����x�l	n)��Ps�a熔&r��`��9Y��7��Xr���FV,��s;hp_A��"�ry��\�+�]a<ԡ� ��d8AH?y��}�S:*�&֎(,�b�������!0O+�"��e�p�ˤC�J�N��o���ƙ@�-���/:�����t+",Ո�����u,�f�U�t	��j*�t),@,1K���b�`ơ��K���-�s0͏��=g�muГy��ݢ� �5%����@<��I�ʽ�e}�Z������y6Ԙ��)?�a%]J���).�3��_oC�s�B?�^�9\�,�c��$�jm<��O:��;R��`A=M�#����v��ǧ��W��e:��&�Rٲe��Z�(J����������dt�"x_$�Kp�;H��|:`��|."&�[�R[4,>�i<�o3ru�=�%+�aܟ0���w�6 ^s�?��sw*�����$�N�#���85� jh����5����/��~v�:xHֳ�o�#.2a��8����I;��rvc$�o��;?q��+\M	q~l&Up~uY���Gxӊ>���!<y��k%f��&��u�gi���T���X}�jQ=i"+J��̩B`��Ż�(|ف��~&�I�#����CW���B�Uc�V̸�i/9��n]D�����&��~:��l���%/}2Q9-�p�+$�S\�G��5��=�x�|����� >�p/��߫��i J\52�tr��^� �	@��@��n5Ң��fDMd�6G��-'L����៎��&2ūs�Pr/R�!^A��aִ������-p�6*,sX��� W:��:.�35,��y�=�s�;�k��	�|p�y��(	8�W�9U�<���8�Ղ8�
���n�<]���aB㊸1*�����?��dƲ��fG!~	�ԫģ��P�U~��z�3���&�>�E���e��	�����@��x�I�#2�l磸�E����N��?v��B���*_����ϳ?��l�̒Q�I�QO)��<� x
�cLXm� ��7�=�>��kӍ���h!8��%6Ӆ���s�>�w%qnqv���4�lf�{\��7c��bhWx����U!��Y��.����/��L�s8��)k�:;������O�&̓ �Ț�Q�D�g��i[\1�W��^�G��d
띺�Z��vev9#n�~&_��[��@c'�n1�$3�)��v�������(ñ������W�<��D��e�8zB�y�~���A���0�
#0��zϥԭ�m��7c��ńF����L���h�~�z2ѻ� ���s���D<���n�}���%��Fs���$m�n����c�(؋�Yb�<��E������$$�W<G��d�Xv��6ɷN��X��P+���Jf;�u&�Qͯ1����~�
�f|E�9��:�2��{#bs�l܄��Y��2;;؜����:�.L*�����݃:Fo�x#̧̆&�K�/f@��P�)N�Ճ\	�x���J��u�qi�p;h�6�(��z}'�*�|.ܶ�yDQ���/<��lEh=����
%mq�9ݩ&m�z�XM�}�dқc,��`�Vf6�+�1��� [�\���/�ʠ5�v?��Hr7�W=��e�E�^([M��x�