XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����N��A�x��*xy�o;��/	�?)3�1$�X���`�Fl��k�����y�L]ݟ��\�,_J�c�B��a�zM�X�5��`�<��7[g��S����B��W�p�6�Xt�9�R�E��[2A{$zY�t���vqe�,uh�
;���_�,���t
[�;��Ȼ�}��^Ias0[�*Uu�;�������N����Y�+�#F �WAY�J�!�5���D�=��D��H(�/�؋0-bo�'U��Zd��n JD)��*�Ȳ�y�p�j>�$�����o�I� �p	�A�J�Yj��/n���l
�����~��N��
�5���|��y<>�Y<�.0ld|`w֕��˫��M!X�z%�[u���O�R���지���}�'��/I�f��B���r{����%���$��3d����,?p�я��*���3%��{#'��xSR�Ѭk���^IoJ��W�#�0vF״AA�p۲��o�=[)��-���W:�a�J�>�[��H�|o2�pzWQ�A��o% 6�t�t�u<�ʱؑ�7Gݜ�̝X=M�j��uF;}f'�\��N�T��o^E�&�zH��`�W=f�ZJ���8@���0����Ɏ�Tz��9�c���ٍv���3�������� �z���t�3�˖��{�cP�\���`��6�@Өs��N�b�6�<����k�k.��~m���&����/_fP�f$�2�W��V�8��, �M���Z�M̹��wXlxVHYEB    3b09     f80/��9�>U����v��7��/B}q|�g�]#�1]-�w5�ed�Mˑ#�db�33t/��;�Q�%!e�za Z�f�����%! ��V�3�D�S��}*&V�mvש@4\ܗ���Ky�S��#�%_[��Q�gq��l�k:ؔ>H�KJO��.�儘CcD�Ryd
�"HǪµ���]�P����M�O?�]��$�H������u"䄞5��Kp�y�|<j�n�x,1��r���U�u5>�W���_E8CI�N�-�����*I�����A�(�2����,�>)�E��|�Tֳ�&8|T$��	�\���_K���d
�b�H�0���S�EP��L8�ԑv�ߍkc��[�? ӻ�h�7�bҔ����-!e�AĠ�E�?�n��C���ՠ�z�gٵ]*�%&"d�gB3E����L��G�����X�I�W�HRsNQ�����P��32VW*xyP<���Sc�C�oH�,��R0�I�����m�oS�LpZB���~��9�pH`51�Ă{�-J�%�g��
,�
�PCǥ�*������i����5ݙ�w?��4+^��7�v���L��3��ɵ�Wg�h^81�R��t"��v���9����^���L&��j,�d�&a�꣰ý�jyz��=��7G�t!��A ��% k*&���_	qFiC�+�H`�������+�oLLD��6��-�司N���IGw�3̆
������G�]�ʉBd��3��	Rp�����Q����êX6�9,�����.�Q-Vtܧ|5A_)�G�x�=���"v6�	c'U�s�n��`�A�d��J�5��譅3[m���E�x"$�t��\f�t�u�ou��ʬ�*���-�@�$��7�?�&I�h�S+=��bA9��BK��TN6�uѫ���(���I5"�����Y� j���z�2V��&�{����¾ϸha���Gj�>!KD��~،Y/�!�P+{����ᒊ8
����D���p�;5�V]�9_��#����&�xM��B�8�0a�ƍ��ш���)���?��3�=�_�H�.w�YWg�pb�B�����Y)�ϯ��,Ҭ8�'�z��N=t�a�]�T��%rH��_.n�	�\��w��T�j�(B	O�������6eO$6Iq�W��x����׎re�o��SY��s��de��,`Ơcr�|�����De]�q&��Q��DE(o]��'Fd`r����i�I
u����T��a�w2�?�W����ъ����g7�{��&7�	w�P^�i����~k`����Nbr�JK�n����:�p�x$8lS�1�ڢ���Ʋ�<�:[�����ُĄ/����*���\W���b����`�4 ox�R�l̩Ea��A͚1�E�_M���@Y�e�H�������[z�H�K��k�rjm�z@o��0�󒫃6ľgc[����yY���~[�o�a�LX��8J���a�\_~�};�*L{Е��,c�]=����(�9�h*��YT��`�#Fo�k�	t�#��.� ���\t��^�+��"��E�Sl�&52�M"���=#��#K�$�Q���"!�Q��r��}�RXJp���]�Ep�ݚ��E�ڙ�hŌj�+��o��뜩j1��`Z�'I[k�\ WUM7'�h�=��צA��,���JB�˜#[�)=���v渆��%����r���ȱ��@}�&�!�����i�,5�_>F�u��sC�辇C�D>� ���p�2��D��I�F?��.Dv)�M\�ڀ_X�W+\¶�,l(J�ض�r=+�˸� (͗q[
Y_�5����J�S��e�_lt�F���y���F��N�|I�"��%�o�>{�/�J�z�쟰Q��	�������`�^:��
�'Ly��Rһ�AQ�N�p��|r!��w4�
�K�)C	���^��L��X�#8z���1���';`�h�~Z; JS��(i ߉����u)I_��T�&��[t�0����}M�S�T]��{ ��$I�Ģ�(�{@��q�̂�!OO�pf*��v��_?��?*<�a��T�ѓl(�&~��`���c���O._��#�j5��(n�瞉^�8k_\���&�6�o�����{[���+���bp]��b��@X?��Y��e��0@�F�R2D}s�8k'~a	y�v��\i��R�*���vs<q��z�u�$AW����ҡ�������r����}*�ɢ-���:�w:�0�(�\_��$)�7���&� �(@"$>����1�y庸jjŢX߮��KY�_����HCJ�Y+�4�ފ�fd}L��&X���}JK��|mio���LTB����� >�`AS�Vp�Y_�v��6�=�����J��oc�j�!���i���Qd������ ��hכ�(5��wK�����C�k�4c�������$X�9�$iMK�ɨ�k�P��Ԧe����.͙`X��/��Ne] ��'��$��$��lQ�3�J��L����2�p���A">�F����	/�OT�4��"9d]K�	v�V��x��Yj
�ɋ�S�h-�l&\q�;|4�+�;O�2e�z/� �r~��[�GY7�l4,Ȳ�H�)��{m��V|z�U~X}�n,%��Jɨ"�Z3��t��]U�VAkt�%�������k���Ե�qf�]q][b�p`�}��(�8�cEd�e���=���`-�iv͜���yw�a�����-&b/P��|Ǫ<����'0'�ަ	M��*iuܔ-���4In"��#�br����K�V�`[�)�O�3{L���Yv�G4�s�C�H��U1��Jl���e*,g���߭�G�iҼ�2�z'��`��t�b�%�=�M�/�BY�������	t~����jI�q2e��SE����yn+�[$w�[�g���ږ����]κ� ��+N���ۚ3XN�c*O>���K^�e����J���xh;��4 ��,�C���ؓ�$X�b�!:(t��*�*���m��g�����n��c>�`�ϭ�y߮�<`�:g �5�5��]�e�\{�7ۂY���� B8@l��=2���t�sn�@q�K�B�_)}p�mR^�l��j��ߵ���%ln��J�.������zr�i��j�����&�/�+Db �e��b���.�*Y������ ���q��)+AQ�\U��˼�,WnT%#e"j�LVN5���d]`:�,����Rx'<�L��|�H��Į�]�n��2N��N��r�rH%1�j��>{j�N(���%#�XX
�f�3(ȡ]���}�\`y�m��H��C6%F�Sv�s���A�Ue�����W�? ]nH�Pi����K��S1ܜ�iS/���!?��((�-E|��:����JY)vZB3>�� w��A-F�X�2;�sVS�)�_͊p�������b�oc�NT>ØW-�P�:t�M�X0��Z������M�p'�&6B�4���U�O�е����r}�N���<�L��;��M��oy<Ӄ�D�.Z��;����t�
�ى6����M�+?k`Vp#�]
����:X�P���Ll�!w�h�� �]���:�I��=�Z�Ld/����,a�![׼���Rqf<���A����ׁ��>�}jO
����P�W"�bgè�� �R/Κ��Zfr���],F$��h������>k%����o�������>:�-�6���C����G[9G�9�g���73��w�P�{�Y�+�������*��g������(�=HX�����]	�����qg3���%0^0�����]о
(�7�o:�Ml�N�ϋi\��E�1j B|_[.c�q[h�!/��i4���H}�