XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��GB,R�9�������%&�_�t 9Z�t'��$�d�͒���ك�5�dV]�tذA����V����a<�T�<���h����	����)3y�0ϫ�4���H�^��ԉ�>����* EX_F}�脹�)����߲�ǚ�z��R�����=������]�v��T}+�zPW\b6����Tr��~�4#.��YT'�^ڳU+���b��WM*9v��gN�eo�Y#��g��z�ي��`��rY	�F�c���+��+��e�`yg���[�?���5=�j"��gѐS����w&0K�w��$�20��c\2ϐ7�GI��)����*j�4���ja�Ņӆ�C�?!��jKث�w�:��/|�Ł��֗����x ��f�=p_��RsR����
խ�䊕��U=�͏��rF�7������f��U(�^^�=�T��`����QK<Y������ыr����R�.d��g�X�3j�ELy&���tbx�W�¦>���?@�y'� Vb�վ����/���bt�uL7��vJ���[ be��^Y���)EK?��:o�0���aZ��RG�$bQ�64֤'��:o}���/_Q=�C-�b�]dV��>�"�h����+���|b8���2���@��@�e�`<.+��B��r9z//ތ��G~��XK�v�����	����i�[�l#��Oʎ��g��7�P�f}�$`B�؍̮�j"lB`��;����5���O�XlxVHYEB    3fdc    1160�՗��]<���|mSR�ˠܑZ�`%Bxc����~k_��N{%��z'f������UQ�>�3������	*>��.����o1O���Jp��'�a� U0E�_�)ݥ�<��-�,Q2�<�V~)��K�bN)le�����Ǿ ����j�_�@2	��Wݪ0^I+�j1p^�K+�����>�C%��E%�7�&�kwNzU�2tH<#Γ�����H�8�Sk���t�EQ��5Ž�Y/���i��P<�W ��L]����S\oǍ?����ơ췘R�T���ч��7��1��7Kױb�s��R�E������
{ErK�֧���"g�����'vz+���xu��E��3
��U��v2$�X2g\��gx|�j�]���S�S\�J-Q��Kk-'�������� !��G��[nAl�Ҍ��7K�n��Sj�����7�B񴥷�JL�FC�c����BVc��B5g���=�ˬi���e��
�P<�׭ن�Pò�@Q����ѩ�bH�[�ܕ��j�k�&_{�x*
x�#M�U����մ6@-�{i�i���ɖ:���tʏk����,F�����/�$#v��FG�x�?��~�xl�t
�ݽ�
C�Ҏ��v��S���~ �j���;7�ޕ��2J�����a� ����֕8H9rV�]RnѠ�D��7�]��!�+=�,�1'VV$��=�h���}K�$���`�N�,>�� E�5�®��Q��э򫫽����Ջ�C�UQU��"{�D�T�v?�mdA�f��EՌ[�Ht3C�aÈ��n �lQ u��N>�-z!�D.��T�1�J+��v3�M��j�[{��wo�,�����ϼ5V��i�����֣��`��B�h��`=f��*�R�z6_p�&`��`�L*����!�`���tgOC��'UjHn����%[S+G�0�"�i�o���xP��mJr�лH���VZj��iҖ�=;I��}'��.�Fi���]����9�A��E�`׵��F�^����6�#�r!t�TB�cD��+�IÍ1�f�.�v2�M	�EG���]�YV���E@/{�O�J0� �0Ē��Aɹ��5ū�Ns��	�`=s�'.�*4�ߞ®��u������=+lĮ���w��u�\���Ģ��g��#��|ۈ�?K�9.w��4c\�s�U�f��$��cU�+���3��0dFQ�*�~q��4�,Kz�3P��j��H��jr��[z������ety��K�"�;�9��_#D�cPG�����V\Hߝ���M<���џ	��gTP振H����=1���El��Y�ٽ9��]��֨>�$���uF�Vնq�Ѩ@�,9��%�vo䟜���3���h���Mx� ��Ծ﷉����oa�9���.����o��iFk�K���\�}.�N����8/ZS�M�r��`)�!���������Z\��b��H�����\G���Kuh�D2��)P"Q��2(o�4Lk�r��s��5�15e2AhI+^��\I��$1���=Xc15�%�?�
��i�אe�u��<����Y����acN�x��3��g��4Դ�����ғ�&����z�W��M�*�;h� ��C<^�M�?[��Uy��\6'�?Ǹ�t�~�2�(�2�Pv���n���ri�&�C�. Z�&%�L����]u*�!CR�˝H8s�В�^OMY�ד��o�V-y�d��gq|'�öV~x���T&U�uy;V&��̽��^q��lY{�	X�ҟ�����e�Dg�$�����G���o7y�#�����*���z3y��u�&���%����	�Pn����)7���dS�,;ӌ�o�ڥO�޸,�D��Ud��{S3�Bx�k�!|�	��1��_�?�M7��Թ�O�w�{�h?}�	����c���sc�P��y��D�+� ����C1r�=���G�V��9��S<O�bn�FcZ2�Ju��cW4����Ӡ6Q�S	�H[�k�5��,���k_����ҁ9��<�b�֌A��N�SsHF��{�G���o'.?!5�����ׯ	��J����Ssm]��Yej��-��?m��Ā��-hxkx.F��P�j�\6����ֽ`�c��	������M�7ث.��!9�Zho͓�����T_j|f��4AȾI�K{�_I�ē�y- �t}ŉ�B��;�`\��*:�vu�c�L���I���$:W�����Im��>NޚM��:5��LŮ�)��&�Å�l$I!g���W�	]����f�NH�/C����Zd3�LG��	�q����ꛯ���k�sH6!w�V2w�5q�_����ns(�e=4(��Pq$�`�%�fZ?�_?:�:�;�^��@_�@ZD�_H]�)[?�erm���w��fW}r���H{l��B	��ԧXL�	t)7�U[����e���2���rs���f8u�������/OW�+�k=��e�;����&ﾧ@#�d����{	R�.��tt�H�S�G�v<�š�paЇ]�e�Pz�EvT��� ]��6��%�a�{G�7X�����7�o�:5�o ~��s��
��=r�{f��$�	v��DK>I�,�Ω�CE�����e������An�f��
����O {2 ݱ��NIaؤ6��\n=��ú��k�q��z�{%����@���c<`ty���<T1F��1@|&��h����FC��a��o.�!|����ߵ�Dey:RQ�y#����kd�,h�^�!	�߅׼/���8�l?����c��VƩ�(ă�j�#;���Q�8�͋�l��
))�d7����#�чs�_�N9�#e����_t�H;;�sHn{t�ͥ^���.�܉s��j�0�1�:��b��������VO��ua-�f���%�7�pO�wn������Rl��x6�c���81��
*���eM�0tW���gpGl�?^�ܻ�R,<��[��@�3gR*=�G`z��ug�j�����`�u��)����9������_-�FD	1�-���g��g��-R\��i�|���'�%2�$�̔�_�$�¹#���}m�g�p�Hp�N�B��Ş��l��8r$?��9n5�w�v�z��(j¨�+B��z���i����zzVf�(B}����\����k]��C�M?u�vD�%[gK
�l�|Z���+(=�h��p���#��Mc]vecB��pK鴘�삨F�u�`*�����^��%b����oqh��<�}+�����´K5���U�p6,�����ި�~�"�;�;��d��m����a��r�;�R�	�5�]���R��qɰ���j�7Ju�~�y?�a,��^�54�It�ط��
����^ć�n�U������L4(����ZX�z��W��$oJ� ��]�����T�dKK1��i(�h.��O`��HRd���6+�W���1`�/uDa��蟼�`����5�m����?���:�C��^l��2!�?wT�T��cz?�*1��@���a�����pP�AK>#�/GMos����%=~g�.��$N��g���|O�$�K��/i�"8�	@H9v�%k��j�=�Kj45B��ƭ��U@�������<9#.!��"���L���i�+��#TN�(g%�;� ��Q��7`Aĝ�z����u�xg?Y��拺��ʪW"_{O(��b�d:m��#��+�& xN���(��gR�%������ig8e1U�O�?���ѵZ�8��~�j�%F�
wI��mPw��ԉ��G���Q�tu�f?�i����g�Z=�_}�}e�
ҽ�-�SNl��ZRূ�	Lt6d}����z�S���c�gW���(�:ȑr"���K�JӇ�t��؟���202�WIf�$�(�̿@�O��3����+����B<{ibf���y,Rݸ�e#m��6��� ���
�ѧ�U�$�n^F��9A�+��BZ�vcCO-�C��$���nO�������P&������A&AZdԣ���ނ�c>��5��k���7���{����	|�������~�a���|� O�l��+$j{����Zi0���Y�d$��fZ9���t�_�e|���%�-��,}����)� 5I��HqiCN �����u܃e�F�.�6�*uE$=sL�"ݞ�v�����G�v�{��Dĝ��QE�_A��	C���Dl�9�]�i�����2���.�o$�!�y�uN����z1����;+��<�qXW?�Q*����K����C1x�2&b	������ODM��KN����:�c�نg���