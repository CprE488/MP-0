XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I0QKe�61�w�}K����SF>B	V���;1�p��;�T�l�9��ǘ�43���w�G�F]i���ȧ�=�e��I>6�k�-C��f#�#̽���iި-:��,r#�i�+y�՘�lОU�nf�|>iE��J���/���Ƈ$��v�`��q.ݪ��[kD"d��<����!]��ԡE�܇`o�E�䭅J^���zҞ#��D�E3U�]��}�jY��o���O����Bq���g/��9������6'��;O��r�O��26������߹^�h��}����݋�P#0���t��湟4W��-�f���KE|0�!���LΤ�|����✠���
��:\3#� X_�<_�*>�J�)윀�S�+�p�GK�O��u��jY��_��i�v{��'[t\��\��dH�Q��׾M��1�z����K4h���޴�I�h^�L	�pi7��j5$���
���5�����f2�4�W@x	�����+�}1�$�a`�A�m�w�b�j��|��de&�aqe��FO�k�ؗ����E�>.�������dg�S�u*�����x�*�Q���[�s��1z�����)�'��~�]���<����mQ��ꫤ7�6`P5�em�����/s��Vx���'B+�׉��k�fڄZo�D|C�u^G�GEǧa�S=�~����
�").m��f�uI�i][?�l�E���

;�g�n�X�BO9�j`$ِ+��(�XlxVHYEB    b3c6    25b0��j�����7���,}P5t� �L[�G�%ri�Xo 
D��R�z+|K]񾋗��:�-v3�����A=Q�/��.�-{�`�fy�4�����<�Fn�+4e)
�CP��ElI"�6K�K/r�mŹ?=WSmO�����2Y���0�o['���vM�6�����}k������]�(.~�w��A���Q���*�d�@J٣�KSf+�a�,pQ׾GX��.���8bw�6V�1���$� M�-����jJ\^c�$G���;��0�!���u��#@b�+�H	��ETU1��k�h���ꔻC)����r��f���f�@³�S�)	$��y�lH�Qˮ
d���\��z��U�"s~]<��L,�C�:�	�@$^��⥾�/W�O��P�zr����lu�m>�j�;f�~�����R��0�V_���%��!�&n83!�������(���g3|������u�E�����}���?q���n �s�Y�$�͠3O�aSjK4k5�99k��M�`(�s�@M��J���&bQ)h5����i�����'�VA��o��tM�X�iQ��Ҽ?*)ib���x"�q�h����L)���>�M�F�Lc���cyϺ||&|��y���=��������\.A��Ҷ���	��}+"�i�kʂ���7��:3���Q�ɜ>j����}Q�����Z��'�yl̉V��Л�����(軔�<�B�,��s�)İ��G!�׵+�ꥬ�K�WS�П�&>�l�ѷ���Yo^st��X�a)��[�mrj���G���i�I��S�QS��ʛ�b��m�í���\�G#?x��>ƥ��b��C(��l��S�黭C*��j:��p`�΋x�c_�`Z_=۠�,/�<Ds�'g�x\P�����k� m��N�`��t,�-`���%���$Gi/�����L;��%�[�elFU�m�����d��*S����!��ͪQ0��!b��	���e���bY�2���%F�39��4IW����!�zfz^�{�raPj���vj����v*�+)�G؉�0:8e�-���e7���;��؛o~Y�[~z:b����n~�/�B��P��n��Tf3̡F�8ޒ�������hGYIP���X���~%,������[G�7���{��7���G9�����H�>���g��͟h0ʃ*����A���p���\�x4���C�M�G�����$��|v��" g�`U�V�|jVPZ�J�aK+ßL`i{N�zRψ%�0�Jd��0��>�Ζ2P�3�"RA�3-�����e{�T�9�\nJ�X��W	�:#=qo���q�i��w�z�BNI�6�FE�I?p�*};$i'�r����L�I��gzDDSe*{݈��/���|�������8�:�GҒ��%ަ�M�J�0��i���n¨�XQ��,�Q��گ��rgl|�H��{p�r�!%߄t��,	4�����k��E%VE��|�uבx����uF`���X�O0p�˿1�'5C�ʈ��?ߢ���bt9gn�����Z�<�e�uJ5=�r��ҮN��Z�9��d�IAq��V�
�Z.�_3��m���L�I��o��6��/ۣL~ڏ
3/��vɊ�j�$�� �EqVLy{F�R���'�Q�Ҳ���j|���F��/�nC���]�)2H������29.�LA�d3g�y��a۝r��H=|�/��y�y#Ç~h���� ��D�ӷ�(5��bae������b�.�����0ƺ��;¾�4v�_��5��
����H:S��F���ꙇ��T�z�<�k1��I�e�$�=���[7�W���>���<��&�N/:�W?��S6���\1`=���Hs0ִ<��$��.��p��cVnp� Ǩ+4E6�T��4.{%ڔ��s���t�]�LKM���Z`d��u�VwS�\��>�r+�c�-8C�9�_M��r��ͧˌR�z11h��D8��������\z�46�B��]����Y-�"Y&�+�I�=��3I>\��m��v����
��a��!�L�36�/vF&��ȏ-W&�ů/�FOT\&�w�ADu�Rإ�K�>�^O����H��A� ^H�g'��F1�RiS�Wو8�;�r���5"}R��ÓD�%����Uk���_jh<*��UW��OgͮVPM�4�8�Y ��;�Ozaiz p�n���Rm"y������Y�����ǆ����{�Q���d��>lp͍��)<���i�%�T}�?*��*ӹZXI�(���q���A--�0��a9�&o�Y'�q����qM~��>e&W�ҹ�0|��c'|Ya �*|�)�]߳Í" ��U~Fr�� �-;�U����P�w�_�)B/����n�~��K���G�?�ñNw�N Z}�KWB�~�Z�����OC�z�����(.��Sj�a�g��L��G�Ꮹ)��C���i���-�9@��_�jѡ@|EK�W�b���Z'v��'�V�K�U�L1@�=����� ��A��W���C��k��I��	�e��Н����r"A.�R�4��@O&J��˚D��}��}���v�������G��a8�͋ � ��/���8�`X����YAdh��Dv�lT��'v����v�ɥ�����2v�؛\ɽ�Ş��o��I�q��)g6h���0I J7�����(� �ll�%�gm����J >��x߶����5C�5����>�aw	�������;!x�M�.�.*�\�Yj�|7��>O�Y28އw��4ي�0���t��;_��W��Qn�!���)/��:uy�Q����1�6@K��ނqz�S��a϶{]���=����&����U>�uXڠD�^f���бjV�a���ƃ���j%Ou=1���O�ܼ�3�'/1"�����@\�`��I��Z�:ߏY��io��?TIi3<�:�q�vi���G\�c;�:�E79T�Ɉ&&��7�� �����(E��!�-h��<�Y��\�_ڡ��$��Q�c2�b(�ōðBux��S�p�&�O�F�(�Qr\&���?����#VP�-^�PH4@V�ȠK���������5���S @�p��y6Yu���ط�گg:T��%�E���^�EO�3�!���j�A�[�-��ÍHs�>rNp&?FT=g�(��Uz���lz���H���=����T�|���R ����'�7����5������n���Sx��|5�^�r�L����d���'xv�f5ge��h�n�{�9'5:�E��w�vR���BEL6`:i�)��f�H�ĥ��E��:������l�灱	��2�����~xL7J��sB~Cܤn���]�V[}l�³M�:�����9����P�W�O��B�@`���Y��$�Di7Ԅ`���i�Z� ��͛���f�ן���A<23�|I�TO��x��K���CEb�l2!��~0ʖ~B	���8�E������P������J����Y���L"�4���?\���a�A��	V�LA�h]�Ue��7�hTA	�|���*້���sDo�rݩba|��/
�j���M0��k�o�y�I���p�K&c���7������{����BrjL�/3��a0��L��|4�ؚMҸ�{�[���������t�G���C��c����ŭyݾ}�Q�#�HQ�{'X`�����WL�9�������T{���T��Hx�ǈ���evR�@��SS�{�����RE��F*�&wIw��_�P匋�:�C�>�G1��ī;c��ɜql�.��B�v�Hq~�$_H����<6�p|��1F3!>ԩx��˼���'��)5��;��(?��W�x�%[��wv���5���t��� A�j�f�q���z�l�ڐG�[�W0�ت5l�x���5�V�f�<'���� ��ތR��Dp�����(�����!Z9�#�
ZwY�-;�d��!�	{�	)�8��IQk�G����P���Z�ك�_�|u�r�P�.Y�O��d��<d�p��9ȿ=�hM������W����ǉ���F3�d�f���1�����������-��)^��4b<[ي�m� ����#'ȥ�`�
�A�_A���8��V.��C�f�;Ͼֱ��>�sb&=r'�D����2G����9��Q�6���b9��VF��"�V�`��]���q�D}�K���2����+é<칶���I,4nBK���Y�Y=AsTMX��ǒ�u�kjb�Tk\�& N�f(ң,_0��ʃ��{J��],�}ǄC��Q�o%į��?��<��$=�"�pj+��LV>]�$��C�t9+v��*���՟�~���,�� �q\�
t:vG�&��~��SUP��0)�~J�\��vvח�|�KS6߭���#�E��
�}i�^O��-��WzK��V�%�'�ZK+䯔�;<�x�`�i��%�V�H�� �ŧu��2[m)r�mpS���F��T��ȜB��WwѢ��y���b����MGr�Ҍ�Uɒ�npqf/x�fE��O�D�����3���}����6��wM.Wk����\[�1�2���e��&��'����)��/���uhROoo�uZtY���j%��I��F��8�$u����õ�7�=w�~������ǥs�
�X"=f�M� �k���D�o�̻�SmG�&�A�2�/�K�Nl��R�}�=�D�ֻ`+�9��x-����W:����c��l�����P�C����\�,��96Tp^퇓<�3�<`� �)�l�ةp�������+�̧_n�W�T��ɲ ��0һ͇� 7b &���hs2F�e��"fm���U��".��R)�`�>K��?`|_�$э��5۫I�}M�AN�F����M+�d!��.�p~e�1]��)b���?4���#���B_��nF�'��|F�-aq��y�����G�Ub�e\)����Ǻ>��F��R��Xy�g�=�Eoo����/���	�l�V�����l�r'�h�G�}�j�Ω��s�}��đG�+5�L	��o�"+NR��{�q�g	���"FR�6�"m��/�$�����y�T��!�;���X-�:�;�%�(�/�E�7���}���F���"�
��yE ��&�x��O��~�=��rܠ�h�
�c�$z��<�	h��ϲ'��PO�j]-՘-i�m)8u�C�Ҳ����F2���%��y������e��*V�U/]�翖H*�]����.C:���m�j�N#��
���v	Q���x�5 !X
������K���$~�s@bh��ή:��:%���F�dH��Z���ßp��5���v<E�"X��ۨ�����!��o��#rnD�͐e5�´�h��,�>Tқ�>O0v�^瞑�eTȴ�CĚ�"�� �*����Bnz��B�~$D�($�����+sZ�k��3a�LD�]���)0XC����!&�$�á�b0�}Ĵ��U��ܽ��们Q�YN���s�g����k� Q9����1I�  ��Bn��#\����H��
 V��iz�-6D�+��#����ć����1��$Y��㴭�!�z�Y�o�]��n]�w�aLqd)߆)o�<@�rH������Y@��#���f``Bzw^ u%��_��R���"<Q�>��X�I�������^.$
������{@sd� 3~����J-��\O?��Rua�h.�m�����B�6yE/����h��o�ىJ��~LS������;�=J���Px�h��a�2 w��t��0���'lԌ?�����|�z��y.]��l�]2T{[���M���;�p$A%V�L�1�@�g���g���y�!�5P"�
atE\�Kc��}#T����j���[5�c�*��k�		
�.��Aֱ��ǩ��!�0IT�ad��;is��H ��k��J�g��[���α�y,��c�!B�Q�O�I�3=����"�Μ/�%�[�98k��uK��ї��-n�|׆{c����(��a]�{ ���%L? �U�/�˱�Q�DBZ;��,00��PxܗL��凛1�1M~�x��8Yl��N�Q�f�_��ΐ(�-���v�S>2����s:O�
u4Ds��VdQI'�*�òD�e��b�9a��P����'��3��B�c
 Q����JO�9o��fr�[LI+�rp%���k�蕨��57 �����hƃ�w��z��f�$W�`�����i[�:-�4�"�>��b�-���O���q�͡���E��1�"sz�����yo�h3�Iw�Z��M�������م� y{���T'���u���d�'G^]���g�j{�ȓ^-e��#�6n�:�����5�o'����=����r"q1�_/o�7,ˀ?��xl�� �)����B���!�q�˴.c���Y�x�E�M㘷̟�^�D� �W!_dh)^�+E�5%(�D ��
�0�Q�;�ǇR(Y�Ȩv[�+YU�p�ƪ��~��s$vh��Ό��Ry�< 7p��WCDR%�8y¸�)ܖ2N���3s�G���/@0|f(�#�k��.b,w*��w��hyn��ٹJiV9ڎ����	��Ij�{[_�^��𼌙�D���<���zF�{�����k+�?O>+�V(rN6�������/|V�rK�}�^5/k���ED��hW !gUb��S�6U��{<�������&^�� ��L`�r�a$��.�ԏ���6S} �,�T������AEJ��I�9U�H�SA#j(�����X�A��S��N�`�X*=�����T��̸��\5��AӒߙ�����U���� l53X��2�]͘dtRR��r���2O�LF��J4�rf�Y�ũ,�+���ɓ�J�!���F������Ƀ~u@M�C�s��7�k����&)v��%[Z��k��ί�� s	�(u�c��z?5i�ٗ�A�OuF�>2�K����l���Z,ӻ�/����K�Ex�2����x�cX��|���-d���҅6�� ܁m�d��T�a �����x�kpxvv� {�-�UQ\��N=�5�~6YhCW�Z��}&@moNs�����&;MeiAl�ա�)��n|ۘ�vf�@T�����R<��j8
�P� Q.t2k�\Gg��^�e�}��u uIϺ���p3��oE���'�k���ڜ����NI�CU�����,NLk���wb<A5W��Ae��2O3�uS��r!��Q�&��� �i[N5=]�Z�� �4��i�=Ln�������L�#��+"���s<�x5���&|	������9J�<}5b&f!�-:Y������m����� ��Yȗ��0&
j&B��R�3S�Ko��)���|Jp���Ɵn=$Od���gr�q���e2h�܀6>�
��H�c�=�}�����]<ȓ���}w�t�M�\]V�3bT�4�)[��
ׄ 
в��W�Xܺ���p��DΞ��r���u�G0T�B �r� Te-{�$��_Nid���Aw�:oSd���t�"V8�+�^����b�z�h�ؓ:ltƖ��<��N��A<�Z�o7C��	��dT ӆ����'O�4�r"&I3r+�ٟ����}l�'��7�rv/E�i3MO&�9y�MjV����?�gn����_����G��1G>M���OW��"�1�q�)���q��Oo	��#��o:c�iIBڮ��r�q���LV{!V�9�҃�C��m���O�%�D�$�*�*��6x���G'��&��1-�z�m����yG"ˬ���s��[QS:�@|�s~�t���Y�v�u�B4Rt��������$3�	FB�Pv�RDiG>�P��=^�����	l�p������n�*O@^:�ã�@�Y�D����úg�֖�$��ɺ����-	;4",ɧ��O.�㭞�<�g��%S�{��չ��`K`vd�Gn�_>�XG�
��ۏ�B��K�B�M@Y�"v͑{C������2��y��!�(���\-ރ�_��!�/�׊���;��X���r��Z�u���p�K
���,���#��[^A/���^þ�2М9���cM�j���T��3�X�x�Xk)�T\�M�6��	F b�¬�<%���T�՛Gp.3 ҳX*_̦5��x�P��&�����b���;��k���}D���L}�
�8�-!q�'"�sN�& v��r~���*�9l�j����b������~q6���D�a� 9�f�y��~L�f`.@V�d��������"Ii��~K����x�@��Rh�>����6�U%K�nM�i�/��AN�����<a!~��N��ޙ�]Dd����?�3��{�7��vĒ�O��j|�o�YdؤX�ᣁ Q�=�?��k]&G7���*��3��j_l �KD���y9-�{�P�s;�&U(@��#�83��գ�ķE|̂����3��Ia�#�b�t�%�#�۬�Ԍ 3���Yu�~��>��Dܾ	�w'�kAP�E=
qV�Uiu�ܬܪ����~MGv	�g�	^�V:��yA�8�y�b�ަ£�����,+�Z*����g~�ÕH�S)l!k��߾���0=���yC�����Z��Q�6���9i(=����'QO�w���G?��@���)7�gƙ�+=$�yGЬ�
�%��pU�hD@�. ��U�
B��}�|xX��$yߙ'TJU�b��+@�+6ڿ�fbG�y/����$�֗/��:��� x�B�"g�W����=�Aa�к�|� wMp��O�)���U��g-��4O}`�Q ���e�9�g������p�	!L��X4O�hR��Ն^�"Po��	�*pAmAd_�cͽ�9A���Bc�iA?D_<ib3惢6\�x=A��/����\�NK9{����-�x h�!��q�~f�y� �=<��*R/�����߶`����=�;�%�l�؋&��$�vԉC��]����_�[#G�x���un�a3�p�� vO��sM�G��;m�}��D��F�*1��͞�A+*��X:���-]��`���~5��^�F�M:��I�g���7��Q���2q]�$�2�1%�b�蜴LJo~P��,Ii9�����.�|���_���+Q����+��v�\u�IG��}����!Ȉϧ���S9߹m[>�H�F4�RߊE,{I;]�VϣB�?!�*���Fjw�,�f7#��A�;��߳%?+<P��̌��������	���fM��E���e��-�x��3�c�a>8�7P�*��lc���Gd�1�;���Ե���1p�Gȵ+��$Ŵ���B�q3���@}�/Aj\���>���U�X�L� ��U���Qr�