XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ad�kegl��%�c�J��b��r)�^Ǥ#�r�Hm�≔:;M�mH9�G�C�EH[�. ���X����k���f޵��e������ʧ^`���R��F��D1��2I[����Ԙ;ο�wl:t.4)cަ���Ve;Y+Bd5�X	d��-��-V�1��#YF�= 	���78��JU(m�x������"n���<t�a��Z�q��o�dq��?=8��׺f!`���X4��l��3��x���R�jR�3}����J��T1Q)%K����"�#��.h��y�has2³{�E�e�g!OX����B�������9� ���h��s��|��N"*��1��}��!��dzo�̋>��ѝK�^��(�y��J�s��
 f'	Q���曒���I���mG����;���Z��8q_T���!U]>6a�gɴ�rqF�N���)�L`̍0VP��8	?@U���J����՞��أr��ɧ��#觿�P͟I��q����v��#C��
E3_�'<���;�S�����`����N�I�OLk��y2%m�+�Q�!H애"��L(��`><�s�#!���?�4�Jw��U�<sB7S&�e�����vA�Q���~OX��L43l�Yd��_�L�Q_opg������]Z����+�����NL#ا���9ɋ� 2��˺�ln��4�>~)�h�ll�5@��y&�_����)�-{��.M��d�W�0��
�(��um��� �$U�$1Gy���XlxVHYEB    fa00    2040�U8�{1p���P~y�(�� g_�[ӏ���[K��1B�a,�!T��*M٦+,È�8���j{tR�9��>�H���h�){�z� I�i�~������`�uˤ<����P�L��Z �I�Ux��(��Q��x�\����>�KA�]VLW��{>.!���"&�ٕ�/@0Q6���Q����Ws�XD��	J��N��W�I����7g2�Ԗޗ��8r<�!s��w� �o>�x�*�j���Q�s	�-�(n7	���0}8��>g�nf�,2�[�g��%֑ݕaz/7���C�c?��K������Ju�����67Q���Q���u�!�/zZ2��{*�=	�U��9C �	q��/��߳���X?���XJ�*`u���x�M{�Ы_ ��;��`�˔&��i7�D�ܮ}�^m�W�.���c.��<���{�)��^򲺡rN�|��{:��/�d큽1�N��>~�� U(['g<hi(!l��J}o%:ҫ� ����/d�H�i��o��4 >����"v��!��N�ы�x���E�O��g�Aa�r*j>�o1eď�\�/w�0	���ٟ3��[C�2�y��N���v�=
{��a�d��♢o�a6������8� ��>��R�"p�D�6֔~c��6�1[K0�`�DvMR0�cw�����@�\�r�٘6G6�dzA!�xC1J�����#�P k_�2̵��J�������M*vW[���G�Ur�܎���!�;B�^踡�o��@�RZ�<sH��ŷuj���kn:$�T�	U麁
<�b�1��u����~�I����s�m��;�Xf�$OH��'e�����AB��"ޖ�M;�xC�n�i����HJ�y-�v1��UM�����~q��DB����C���:�|��I����\��Q�$��8a�~}^!/~�K �n��&�E�TV"@��6����;Ѭ;����ǒ1P����,�p���@��>>O�l�$�N��&��ؐT�Qe8<��F^��Y�1������dQ]�.ٟ��KB�F��Sn��h�pbwīq:�#�a<*��w�������Nt��b%h:�U	v�Gs;}@����}�2���> �(J�IwV�� �x*�ɰ:�Z�����=Z��JO��vXk�赠rn�$��o����[T��	�ۏ�֌"���໷�Sd����:�o�~EI��r�9��4��CD(����꒨m�]��6���(L�G.�+b�WC����,>Pe9�/��/����i��#�K-�m�rp/�s����>�/�.��h���L�xt��7��⭀�ZO�`5���+C��BW�,��ލ߰��ْ�ϤJ��ܩAR��w/%(��2�On&����p����w�G��r��Wm{���0`z�f��\�o�UAm�C*��X�<\ct7+�xur'h���:�gA����z����q��c�bo6C+�s�t8������=�:�qR�E�rҡ�+��3=8Z?*�V�ݙ&��+����J�+��)k���Zj���jk8k��&�?.��Gq��~�Ϥ/ԻY�ރW��A���J/0�Zj���*j��a��l�s����4���#����U��~%�6tVk��S� �ۀ��
IPAh<�5ng�}�(m��"d�7&լ�`��/$�n< C�o��j>(Ꞧu�(.jG�T�(��q�M�7��������M�:na�e`�O�&(������H҄@����]��8���b}0�9��a]>=|��7��t�z�;�y}a�"O7� �ι籝��Q
-�[Y4�=�2i��=���� �7��VU(����Z~D9S�	�q��.���R�'ɟ ��܇lbIOwՀ�:�x�?�説-�q�jD���W'�ke�/="w�/�����S�/ �Z",�~�<���xsP�j0_]�{���JI.���K(�e�s�<�k���Y:�R���r1Uu��󡲗Z2���:��k�cĚ�K�������bT�Q]���ˊ�0-~��(��*:��JCN��,5�����pK�������BM[F�J�H��Y0�<����	;:Z�(0V��\�Ύk�7��E������ά`�b'x�3B��9	�v���3w�Ͳ��i��Ok��M95�����^Hj��e6�'�����7��,w�;�������z�
�6e薃�!����s*x����yOG׆p�D��� |�IE�K<��`���ȱO����H�d�5�A��!�=��	b�����a������aq<��n;/�]��4!Q+,�v�����@�qܐ��mє�_A�~8�SI���&�&�M�b����h���x�jŋY3���LQ8;�L{���Zl��!h'T��։X�rXwI��|�d��
ᣉ�m��ک″�
��]]�9V?�������~)���E)L}�>�U�!۾������2��m`%nx2`��:R>�IXg ����}xh��)3��R
�	=;��y�g��� ��4�	`����Q�
6��:Mb�":� �1��=�
u`xnh�޲�4�6�����ur�!�<PQw�D��Q����	�\�9"��0go�5��d}c���~S�*³�ӆ�">+��'Nr�;l���G��e��abmr��)Aje��{�/��(����b��C74{���R��nH�q������V�J�n߳^m>��'Z�r'�O�V�q9��D�<����h�A������bOI���M�+�d�6��$��+|rp�m���2ӡ�j�@"�%w��W(��������{���&%��bz�(lfz�pX���B+&��_nJzPk����t]D�F��uh)S83�F�Ϲw�>����6V���#�-FCMWajkYZ"-n5�FV�0��@��L���	����ݮ��֦���7՟�|�<c�K͇b7�C��=G��-p8�����@$s����\�փ\x��N�&���FK|����LL��hB|�V��ӡ<N?q@���=�D����2��<�͞��Z�ρRH�a��&m,�A?�}����3�ڭZ&y��4#L�:4n�8y���̝Y2�G=Bnl �\/{��S�Oi���')�\{�;_rO%��-��񇚳��
ȿ��8�SG�:8c? ]��ʕ�c٭&{�S�\���
F�ۋW_!YL8�#��ٲ]{|��u<,>���X\][�/Mf
�t�E�]��4�y������9pX�y����˗����ѕ�j2\H&
�d*}ީ�R�[�����Pr���j�p^�����4���D!�!�`�N{UP�z��OG~$)���"):�|03�#��䫟ζ���J��{��A�z����%+
��҇�G�Xq�UY�}�$�bU����%�a������_�7`� �?�Uϔ��{��vWѧ�b�o�X�m<�w�F4��6�R��>��b}�-�9n2 ����B����\m��ey �8��=�)���E��9��5PO��0����,�8(=p%�s�rÜR�Ƭ,C���ֲ[�;��(8�@>���+�pmVT1,��F�j1?�o^S��̞{��Fȱ�H�;N�� rŪ�R���i!�,���!&�׽s���`�[t.D�|�'�.�@B��nA"�WUɴ2;7ۿN�\�5i�wN[*坼z���5F��Xu�8���
ǜ�<�b���Rn�zq�u�k���q⣔-Y3�G��,��x��\���I��1e�j�/���ݙ���8u>��Z-�P�z��,\��ٲ���R|ӘP>:�X�(�f
G�B ��>ty�x)%ѯ���^=�[x�}�Ҿh���Wٽ����B�x3��{����c@+�R�e�x�����U��r���8�0���,<G!n�ǵ�;o�֔{��ʫ��%W�l���@�:���kR�&�S�|T�C~wYQ�<K��p��1�`��@��5�8��a`*��1��`D?x��BDHoЋﶟ\- аp�u�f^g=���
���+7�6Y���uͺ���������U�9܋(yn����Ï�[F+c)&u�������9���z��ˣi�U��y}���J3A�[�]j_��o���e&��#��/@o�,����"(��w�!s�CI�8��Z�iK�n%=ߪ�Gn˄��ɿ����h[yA~��MΦ���|l���%��\̐��m|�gn�c�~��!o�7��&&��1#��O/��g�h��g�,;��@4�֚�c��`�6���pH�b���ײ�#ՔUV~��M�K}Q8�?o���0X��=�����S���RM!]��G/)���V�����`��b�@�CP+�o�O�����j�Z߳�Mm��睊ӡ�Ц�����d�چ��=��F��>�U`��ު�K�NN ��*�ޔ��H%�F���Ff@ՋN,$|�n�u_�.�!�$���Bz��&;n7��]wv�lVϤ�>����[���0����mk�o^�l��5�ꙁtzX��	@R�q	;�3�F��� �f�3+��:���}����|`��󈙗wj���R�3���F��,�kC��O��M�`?| @P�����1�<�&�K?����I-:���άI�FhY��G��>Mj�x�_|�̡U�UL��iܒy5�[FQ�Cz	R���`y�o'��=�Ěf8��.]���k�㼚�`3:�����s�~��U%�P��̣�w�Q5Ol��L��Q��T�wԛ�3TS�>�.D�<���!���+���,R4�F�!�湛�u��ߍ���� zÒ�|E�%I�`�Cj�o��;�'�"黒�i�գ�i8��ʻ���߅��E[G���ph���U�Ȯ�|�ʮ�]Oz�<`Ff��.c�n���w�13>��,���]$*�����uX��q��)��F�z-�	,`��	c:�w�t<����7p*KR@Ce�Li��� $�_��k�l	�2�o��<�.��9�|!�#��y�0[S�52��f��C���@�(F��X�5�nq�?+:�S�0�����R<	��K5�et��2��iH�0����h�'+�gnn��M��p��T����lS �r$ɛ�j��kϝ�r]�]��Ͷ�k�9�:wk���h�i�Ԁb�v��U�
#�vu�ױ܁4;<�i�����+=�i��k�I�!��C6`�뒔�rZ�m��/�#Ή:�p4�C" wU�x`�����V����l���n�A��n�|��mЕ�Ü!�A��Q��VkZ����`�)��}�ѹ�Y�� ���\�0�"��e�1�j�Z��;�}�J�JХ
��z�Y(?x?1�Ů��:�_�K��8B�{!�Sʴ]� �2�<��E�Y?��[E���Z]��E���MK�ϊ�.	A�%�M �����#���4+��B��#��5=�M��sc�W
��MU�9���֨��I�i�Xa������W�<��o�	�x��6F��'��ߪU�ܛVM��+�v�� G̿�A؉�W�7��b�D�Y2�Q*}��g��(2�����SD�Pl�R�[�F*� �q8��P�<��<�EP`�j���~U�(�^i,L- ��u*u?�Y8a�	���������LH � &·��9c��oj&2� �M!�p�7ᔸ� b#a�'�����X��8f��ι ���߱���'���å�2P�Fۏ>yM�Mϙ����o�0K��3�t�i�,d|$G^�X�ڣ���>�}kq�B���@���WQzF��!�*�{wc� .@Qk���� ������+",�J��k�h��A����Xt���.���� ��~��6�[	7�7B��l$�����J&��2g�U��pxk��D�P׃J]
�$�L��G��?�_P.1!�j���m�w������h�>q���z�HY�����x��k�c�x�؃^�+s�H|B���;�;	ks=��c���k�� 3n���bu�7S���CMa�羭���"3��v�[�񣸾)s��&�&��$}�C{�C�
�(gS23����l�����#�����W!�&�I�v��������>5�o��F����.5�Sv�_�dǎ��+�{s3~nfs�����O��u����������p�C%	ufOPv(`�B�'�D�l���ّ<DDX3��ݜ߼�O�N�	�hv�ڊ �EM��vI^�3��4T�#�g��Va͠#�T^���A��C���8���e4[��|��yv�4���y�u�A�ūL�Bb�cN��U
! 
���Á��	d��ɭ]�s���"��᫧o/�4+��i����䓲�����z�-N�`��h�L�^�[�N+�h�����x���]�5L��������ݯ�P/{���4�ԍ��x��G[�U�\�4rY!�9xD����l
��R8=���=� �]�lo���JZ��Q)\�wM��d�� �̟�^��\���hiA�0Jv�:0�--.M.��<Ȩ3��\����$x�웑�U�l��8wC0�b{rM��\�^�S�C�:5ze��Ǟ��)�/s�H�f/��ڃ���@��<lβOY�9���$y
����*�,ٟ.Ϟ���u�*]y�w؊���0��KO�L�U߹�F�"G}�n�����3lR6��e�v�(��y*�t;qA�C;Mر��a0�<C�{Y.�Ħ��&��v�h��h7-]Pu��'6ɚ���1�~��r��AF��4�z�ҷ�f%�C_tn�1Rğ�=EAN2�AY3w��M ����	o�V���26��H�FI��K���QM�UR='4R���-�}A�L�Q]Kj��b�@��=��\B��*s�l��C08nx�F���Ns;�����B�O�V�ʵ��*LT��K���kH�Ԁ�vo�r�ָ#eO+�o��,�JV:1��}f)�H�q��A��\��Y�&���qSl��{��H9�be��]����`�p����3og��&�0���1��s�Q�ml�]p{t�I��5|Lo�?���S��["#�+�P�tQW9e��)�BJe�Xӹp���hr��z���^ܘ������VA?�ik'�¬K�o��+9�<�j�ڿ�x�/W(1������\U��M���	}gv�eK��[$���L������{r-���F�P}Rq�G	<+��y���JxL�>�׵?��1�h�<k�廖�Z�O%"w�=�H�txD��� ���h���=�� e���Z���Ӓ�J�����p��)���� �h]s�o�\H�`ˬ���Vv} 0��+��j�У�VRe ���]/�||�M�������e�nH@x|�5c�o�k�32�������f���?�\&!��J+e�����OW�[�:��y�Y����_jn��%`�띎�ۨb�	�2�]�T�m)O�6�mޥ���gg|�	tC�
1j�,M�ޮ�}k(ߤRR�+��$L��"q���J�}��L��_��O�����8
&�5ւ����)�%���'��J�:g����Fl@y/� �������/͠�k��|���.h���Ut�e=|��YZ�:��*�#r���W�3�e<�<�V�$Lȯ5râm�>
�R)��������%�;<ĴW�
;�xW4LW_O�e�:hq���~�_�Z��ez^P�k�/�XЎn�"�,�!Yd{�� �B��s�=����_aO*��և�Q>*r�Y6G��;�7ō%G;i��q�Ud�N���S���O�}�.7��-2��U6d�7n\I[��`.�6Mf��m���ߧ"KA��WŽ��$y9;a��k"��t� 6s�Q������Pәp�yh	\i���ni�o��
� ���U��L�?���P�EZ�GᢔV��m]ʏ��7J�>e����z쥂�)|�I�2��}9�zx;{��s�G�$M��
#nP) V�p��oU�.�5�]�m��췠 �oK��L|s���mxsA�jS�6o{�e�\Å�Ш�1���ij�9�@�xWb��>��G�<�j���>�<�o�Y�6ph���?�2k���<~.A��ܿ�r���ִn�;�(%o�0b��gS �5�pXlxVHYEB    4f62     b50$I�@+�;����ka#�W����i(Cp��W�Q{m��ƪh�Ŷ��wv���X�f��=>��9�؀��ߧ���Q7�W��7�,��6� ������f"M	��~�U�,�3C ��Alp[P���շ�"�b�%�� �:�`攌��j��J��45�=`�F�FIMn8lp��2E#�k�_�?D�N����!��3=��Pۥ��؄�ar�5��|�2F�u|���q�*��Ly�X
3��Jy�M���h���q��O",dH�6�T4'�x��ef�)!ul��av�v��,�o�X��)�H9��:,�<��hb�S���%��TX���]0>0��8g3�8C�ֳ[i�C�;U����S��im��~?��+�ͽE#�o�I�$�ëx���P��i?�=|�H2 %������K�IZ��});n	洺��D$��w&��6��:T�o�=~[F������$c��p�dQ�Mi��  �b8��d�Zn��!�ۯ�&D���-S�׼=���͐.�Ź�_�t�:�0q,��Q��au	��f��q��e���5�
��2eW%����^g.���n���m}m��I��@�z�=}U�U�s � c�f�G{ǄD�JSӧ	.H���쭦��g�ڿ���� ��8~�{+ݫ��O��= $��(�1u�8�j���l�Ҁ��lY�td|����1�%Z�w�W�uj���Ǝ�+�� V��q�;1@��TE؆X���6A! �̼����R[�ߣ?��s�J���zF_6@�)��ȭ���w^��eyku��ԕp�O��B�����bZ�������/��2!�l�x�8���M8pV�Y�D��c���*� K�C�{ƕ�:�,>�D�<�A�V���N���rI�� �/B!�l��z�?=��bu�<
}&C��.T?�2K�~�}���	Y9d���p`�	�����4�G�C┿�%���ڶp�Kb�"}eȼoln����J:�A)�(��`�U��d?�7�H��.��]t{��[�-��Zn_�ڥ���ѐ�A+{�S:?ujo��%���&��o��5DK@(�x�ȝ�,&���]7���u��� �%�sn�<bd�-�*D�P�F��C�Z�V.ݶN�ȳ���FfY�`��F�#���T�ڇ���]���(�|��7I6ҿ�q�y%?yy����|ڈK^y���| ��b���7�Ӝ6�鈬����܄hyJ[:p�h0<��$Yq����1G����%�v�f�t.��ry���/�n���@v�X/��3�("�#���e�ȴjShʰ
�}�?�_jM�j|�%�~��p!d�{.�f���y�٨���
"L��� �w\�W.f��f}�ު;Ŗ�e1)�a���l��?{װ�Q��́�E��7�t�3��z-w_u/
vĭh��L��s�eD+���iix֎���rl@}��{��&�[s��?kRٗ�����G��_��rTvDݲ�%(�[Vg�Tv������C�agv*V��j4찺=E��Xi4:o�*�2|m�q�s(a+42���d�[��-�:DG������!.t���a��j!d�=X��t�]�w_PrT.�9*U�AeoH]�|qܚݙ���`�IS�^����8-��Y�k`�J�+��e��kR��5�'��?(����@`N�� ��!G`���ϪˎȖ��<�%O*���rB�E�w��r��'�_�j�X�|���Њ!�,�^��\J6|�"��;!b��l;>YC�x�k��=�{���TUi��XU4#Î��Ϡ�)�a���̣o�<�F��_F��u�:�h���'נty8���o&����iX��.j�NIϠ�d��N��p,��j��$=�uɿffB�Z����}:&A;���FU�7�gO��p!�G(�)�3\[+�@���:*gR����V&��I)�̼m��j�.�N._����c�K&N�sj��BTh��J��Jt�?���k8���A[����X�RC�χ�D�dl 媭��=�*2��$+
*=X����s5���?�d�_��������/�<p�Ah򨣡��t�h^�F>�wa���i��ԙ+��;E ޜXCx�Q��.GL�!|�Xȑԡr>�KJ`�m�T'aYn@N�=6�zS��c�"�m�+��J*_ߏ8��#��]u/��8��1���T�Y�k1��=)�t�0<�.�Q���0Cqd庯d5КN{�}G��l����#K��P���d�0
���5	�3z�+���5p�I#0N�qR�_Vݕ"�O��7�n���/r#�[��M�&U�*y����D7��"��i7D�J;�I�,a�]�����*[��U��o�ŜQ�#�c������A	*��c��viL���-�t�����ț�o��f��}M���9��,���wŭ�(�a]�G�������s=�;�CH�6��c�j,ave���H�D}��gb�p�J�-d!��M�iU'`x"��W�1��mN8��Ή�}��������0�[�tj�`�FO;k���Čs��1��qE��0�$�����7`َnS��G�,�+����kA�S���ND�e�u^������
^mǿ~a��6x��E�!
\�ɬ�b���~O��H��V���������b������qg@�5�[H��9���}��2y&b�z����9����S���b����.�=�<�p�#��Ƅ��K�Ӑ���~��?H����my���X���ai�.gykJU����ډ�#����֫��N�C��)V���q��&���W�@��Ԇ_�!7�a�&�f��ԝ@��UfB'U