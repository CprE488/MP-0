XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g����e9`9��^>�5&FFkl�gV1|�WA� ��z���p(~��INŽ�S�A����O�6/��p��\Й��]�x���XEDW����,f�vk%��] �c#����@����Ƈ ~#�ʊl{B��L{h�wr�(�`;��s�>�wڸM:���!���\Xp�^)V4
7L���~�ӎ���A��Hf��j}V��?G�ag��L}��w�7b�۴v������k���v���)����7��ƍ6�NTZ1�����<sD�Uori~��R�x?d�x��a�	,��4���Tr�G�G�>0��#u�"#�Ƚ>�']O�+]��4�Cr�1 �SFb��>6��,ě��T9G�?�c��2��-��k���'���\?��{�|��m�vp�# �|,.m.js���<a�mj<�� �ѹ��&�=�w:{�}�3�گ�ܿmE��&N��Y���9�h�%�񃹍݈yw,���� ��Kn##�D����l�Ψr�%#��s����WƢ��~JK�v2���8��+���<�J7��ܔ [���z�${�;)�X�S��X��"��} {��5nsP�,	>�Ҹ�/�!iE�ݪN��Y%��j��493S�>\���_)-NGhj��=n�1z?��f�ؾ4p��yz|	��R�qYꔦv2�c����a��7���~]Ws�z���+�s����o�c^YV���H4���]N�{�`8��-�ړ88��.x�z�	����I�%�b �XlxVHYEB     f6d     6f0��'D`�-�om��?LV~C�^*LSg�6���� -W�ﰼ������b���R��eJr��\�bz=��CU)���x���=�����m��#��s0m�e��Tj��F��~��'3c�H˞Du��6
P���+�����G(p��-uۄL��_�d�������9܇?�!�f��T�\�n��� Q�5���a��'1���W�r�q�I07�3�P�7F��QG,��k��2���R�i��X�	6|vHlxB���F�M�3��{,�)V�Q��E�1yo��rB��k�6�]�����S��ৣ9K|AA.�B����R� ��}��q���xZ,��;2sΨ��V��|}@�d�w��Жse�V�����0�� ~9�󊍟5q=��O�a1L]��Iu5�K+��aw�� 1�F��&{ t���8�2�I(Ըݐb�b����#��A��U��/�n�]0wv��}���.���Ӆs�#J2�
�KpF=BD[�"�HÞ��:�~a^e�M��J,��f19�����:��bp@�g�IVA8e4U�:�Ũ��=y
��}1ݏ���PES#M,�Iw�k>)O㧣 ��2q�{5�.{��W�4v�`
y��>�e��݀{��?�6'�J4��ǿ�w=i��d�.��A�)����U:`A+8��7rg-��^<.ܼr�2�`rL��KQ�z������h�	[d�gX&�!?���� {��]p�*ݪvF�/s�.�s~�3�P�+��W���͈$p��j3+\`;�=�]4
���Þ��!���Zf�c��R����y�N��Y�>q<��}!r^���ن8���t�7*Ǡ
pj����J����p���R��䪖����+�5_��g���t���C��c����y�q�i�a��)�BE����8$�N������N�G7B���èPED�>m�;�I]:�M2%<\4�^
"��x=)���P&�n̤m���,�R���*�,@���O��#{�}a1n�U	�v����Om�v��+�ć��l@&��1�&,���. p윆|J�8�M>B�F�^Y����~D�
*l4\���.��\�@���b�P�����mŚq%�r��
jN[�;i�4��*<_V�V���=,���ܬ=#�웮z�u��^G]�V$�S&Z�3��l�.����� ��tq���iq78^�(�=@FIt4��^0n��%��2{�޽p\}�x�(�>��&ί̑'��(-��}�e1/�DD�G<0Y�e���/�T�=5�xs��ƭ^��T%zuM���	��5��H��z�6�C�@�������`�\��Y�zlEǬd��$�N�^��G~�ZlpW�f�֨W�l�+OMF��k�5��:WH�����*T��W	 ,�L��d�����"����5]��s��S�4dw���[5���%T�+<��nj}Iռ��1)��C��Ӟ�n���,4Y��%�P���84�ؤ�M
��!C�Hv,lP�*WB�����ǖ�]C%�~��`�Ț@��A.������ǧ����K"�a�'����ja9��
i�o���Ω���6V��o��ѝˋ1'��&ѭ.k5�����ɮ��6���P4��/��C�S';��
���Y`��:�ZNۙ;����бx@ً���زj��o�a�#�c�叐�2z�!�_Uw����Օ�i=�%n@��7W���vz��Z)_�أj�%�"�A#�:n�B���f9�*>�4{�:����f