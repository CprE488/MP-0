XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���XM�H�:]�@�-
���=pY�)�t�9@{�y�
���޻65�84��ޞ�_���φ������Tj��R���)��%���?��?�F:r�h=q��;�fف1�=��ݢ��Ρ]���-`�7��/��k�/�=]��O��;���D�Ms?�y�r��&�nO�{2/e��h:��v<v����U��miS	#j���sS;S]��	\�ą��>'�w�^�4��x\�g����e�����LD�к���;���63�9�뒏^V�5	��z>�����?��ʘ��W3U��������-��(���	ī���Hyg� 7Zo ���
)��6��8�-�p�����6���WT� ���m��:m6�_P�����_�@�H�.�t�E�`��Q� ��>���p�r�d�JU�4����Hٔ)>�bϾ�A�
�J�+���v4�>��w��;�u"s��K��Gz��i$Ce�r�ۅ���i�<sȸY�R�;㹚qt�-��{�L�!�?,PUzD~�L���c=؀
�n/)�����"[� h�έ�V�[��ҺB%cg�Z��߲��&~���C��.��9��rf��|"e�@~�o�gzZ͒�����jN�ʺ�7V!��>�S�r�����#V<���K߷c�I��8�^�![Â��㷭�J�4a��,�8ז�1� ����S;s<����)���
��3f��s��0�;��1um|�y��WKXlxVHYEB    3fdc    1160��KvXV_r���-v{B��a�@%�} �ڕPn�f�fL��6�:�E�iB�n5���cTV��
U�Z	E�B�B��
�,jY1\�#���r瀦��y\�(]�k�ޏ���=s$�SI���Ź��W�ts�b��E;As8{����B�@�/�z��oS�*J���U����qK�Z��T�����~��y�#�m�z�tA�O���R�|p�U�����B	��e��L�m�L�����W#p |�2�D�>��w�b�䌖��e+�N3����d��J���q�F�5�=�Dsm������J��'!?�߀҅��8�R�'
���	BR�}�p�5�4�@�*y�<�m0_�o�!���X2��J3�R�G�����=��3��
sȊ3G%H���Y��8��+=[�w,#�������gW�n�U`��@��0��3�tF�9���G
�Ã'0���lƪ�4��~|Rb��kƜ
D����X+��^6�,������%�~K�I B�^+��P?C�"���(7����w�:�'
វ:���8�T2�,�Ջ_C*���Q�}V�D�^*K����*���[�:�x��睶�X���,�gT��A�b�"���⫽g��B�At��'�_Q�+��س����<���X;�
���T��ʻ�'r��\>ا�T틯	���fh:���6F��t���k�d�b"��.~gs�t�^B�MX.,Tb�y�KNL���ɕ�G���i��N�
�M�R�����(��L�k��:��f9R�yi��T�O�;;��D��"8'9e��`9A/��Bκt@�^���kų�l�R���nF������-����9�����Bl"0|I�ƱN,+]�	Kf	x$>��� V��F�cqVw�P<�l��'qC�q�͂�_Cx���"+G�UM�Y�ph�ze��x��@s'�ۣ����k�x�:�0ĭ#C�@L "S�2��^�K�f~���p�a�	%�ɀ5�lz��gT~�T�0IE|��6�(��`��6 ndW��Q��X"ߪ��Ic�ul���V@��y��27]�>v�7Z�H2��bDE��N���>�4ݿ�b)�Y
���,���O��;�	7F�bz�Y���q:"r�0��upȰq�%v'_gOu�8>Hl�:%��'F�ᛳS�F�%8.���y��7�8���hZh�Uq���>>Y��P؛ʌ�1�-�Q�e�{+��A���eŐ����K�ɱ���	�R@X8����BK �E�v�����%��"����x�p��l��H�`���{\1
 	����T�!*�� ����3GBS�n�ͨ��
8��,!������#�}f���W�h�=_R<I'�ЪnyT��QN�x|��p흸��&�����P煛sm�.��Q֓��w~K����\�T�2q�-c#5B�xh���Dy^�\�a��S�ۜ�޷p�H4�ٖ�-4b1��|yc@(<�q�X(��Yv9����Uy�3p|��p���q<p�OO\ ��;������>�_�*|_�yǄ�uC��c�pƜ�������1�IK��|�,�#�K߆�L�Y��-L��(vfX�M_#�3�Qz<F܌]3�֌��p'����cT?+y����i��f�����j�FR�NS��a��<��*ݶ�f6	��-����ґ!S�������0�l�""���U&26߮�\��Gf�ߘg���3E����y�'À��A'��}%�Ka�޵�YW����knJ�&�F�^��W>ܬ�&s�o��ҍ�d�VJ�����������q�ߔp���&�)��`��M�mR�L
��h��ϔ�]Êz7	l}X2��+̊�=��״��b1T�1������*��kf�I/=:��Ht��*���(�
3���uq�df;�?����9�F�#��,7z�@$��{Ӵ��2�u�c-�p������i��k����!YŸ=^}R���bt��}��o�4]p�W͒9�1�V����&V���ϡ�m
%��/�Z�r,;���a}����yrW�]�����i7C">�9��p	ZX�g��^�"��
G���Pg��@����3���Kt1RM�Y/5v��v�0���7�k6���ٽ5��ŀ�Kz���9J"ٜ���(b%-��kk�u�G�>��ў���W�LC۷U%�رbX]̡�<]>IR/�m|�����n�����^Yh-��n��`���>�XY��#��޿#�r��BtD����c �f��OJޫ���$i�[��:TW���s��@iR������V�A��g��6�_�e��
Rh9��6�#�2		��]~G�N�-��af�#W�������s�~|�o�ǥ��q<G&�L~]Q��vw&�e��%b�]�Aɛ�7�S�J�%�����c���X�7������B���OW�ɵ�,��#�Pl��4�7���G�f$��`>�L�8E���v�o�Pd�Z?
��2��F��i���U52�؛�I\O$�<��ࡖ;06�c	)��/	 ��V�(���!�)>l���v
�ήy[���%#�������4���W�f/2V��-� cD%O֪I��m�w��&,����
*B�H�W�p�]����@� �<��S�Z�M�wf�Ce�����7�*��/_�a�q���t/P������g�pe�{9�t-g�RV���Z^������{X���u9R������ݭ���"��e�"�*��hD�?��#�J4;�X��Ο�<94�y��5���e�����L�n /GM��(*h8�F@��&��S�p���_�>�bKK/�r|�d�p��Y��u�����hcߺ0'�Q�F�r^8V	�]��g�9 ���c�I�^(=�S� I�r0�ܩ��G_��\|�^
�0����G����G�#��'!X��w�M����40 ����9�7$��Tc����`Z{~�V\��E��{"X��n�y�mO�_^���M�u�H�'z�rM��EȡX9#�õ��dMnm������$��v|�K.ޮ��9%�r�(婋��a`�V�H
f�I"2r���p=�&1��Sʃ�����&k�K�Z�y�<�F�	m\w!�{�Zy��*l�������A�Z5�r�㥊�@>�7�u��TM�,�,ߣ�t�K�f��i��d�.O�SE(�l�/t��q�9D���$O��D/[/:��9(<�P׻.H�h�#b�G��A�4�2n�i7'r���H^O�����rW3�� �w�ӄ��j_,!O[��%�#6%�[]s�E��:�-�uAƓ֭ȼ�� ��Ĺ�H�Z��6�%�D��3�"�@�#I�y���6E����s$��sV�8( ;K���Eq^�#�=t�؁e�'d��X:�E֫��t�ؕ� ��v��H�
�s�o��Ð�m�NI���D���O���N���=�)V��<��&�UV���3:{b�%�;����C��F$p��4^�9!�1r��\��Bf��,�+4BT�4����]ǿ���u�p�*�u����p��>/��D���ߪB3��w_�$욁g��%;7P ��4�9�v?+>�J���ݥ�#�<���qաԹ����Wms�O��-;}���$Afk�V�1F�{ (�zI�����\��J�ת�ɦR!{�G\/)���eHEX;��O��9��ٷ= c�6S���O�S�XR%�BUX;�u�p�`��.� �����X�E��w=u
?h��A6��o��xC '��Ne3�E��T��Z��ioų��|m��w�Ю?uԏ�2q�/�e�]�9��m!�OV�kO=���␑Y�&A;L!S�Q�f�:jK��y��ꠛl7��c������f4�.�!A�G���](j�Wռ���'����6&����&4Nص�r���Ke�]_#ߝ�_'W�E��/\��r�c��������dK���(��1��+��n�ɘ�R�G�ѨEz&�#�E�㲟W�?^Sv����Y�	XC�WGͼ�	�rTk��?��b��Þ�9�mݍڮ[a���bb�������xa�G�ɔ�c��t?f$`s���?Ѻ��wVLHH��T�ɸ�r�,2t�� [W:���<A�L)�+kC(��Cp�E�ޝ q����HЃ9���4�Ը�\�@8��:���<>�,L4�#�G����fo���:�Z.�T�o�o�Q?�&��߿�TL;��F0����_�Z���޶��� ���>����"�{lu�ޙ��:�U��NQd�$+^�t�O��=�K0���E��� �U/sN:]�f�F$:�B�}O��e�j