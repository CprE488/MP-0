XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��d�.8�z�lQC��w\�W����=x�м�wmЁ`�
��FXU����/��1�]q?�����me�S�؁���E�/ꇺ�(P��&~���li^D�[�J�ɇ����ս�%�WYX ��Ȣ��ݎ��X�DZw^�7zv��>��U�����o��k�	�q�^�2h����,���"���~������g���Ҁ�ЇAe	J�&�t��׷�e(���v�v�{�%\�h�2�Fz���0H�6_��h6bT�*��4y�g��UF_V_�(e/!���6^�F�jY5d�*٭}��m@(`
��0_�u�n��i3�ʖ��>j�-�M=E/`���dċ�-WF��:��
�u�1�AW5���:ؒ|73�?���0���@j%������ge
�qfr�G2����>E�!��n;v�l:g+HI�0�}��{�� c��o{�+_��o�s?���ජ���Ibpyq�2a9��K�g�{v:<}������yh2��˶�Tד	pC{5o�V�Q��e	_�icX�Q�!F5�ėqC����Z��6���jWxnpQ:��_���۶�-�K���EE�k�kq�n���0z.G�7:��e��_��ȵ�C�I��N"���%+m�@U	��M�r.�fy�}"�:L���0��~al�jm��:�pG�J#�M"*���;:���"G��JFS;����"g;�/$������w�Z��g8'X5�_(���@H����Hj <�c��C�ŷ>c01�ܧ���[�XlxVHYEB    b3c6    25b0"Z�k0�]Vq�Q������ƛ>~��@n!����p�U�	��-����
��A�t�?�~���/ WH��P;<�G�b^��������^��P���L\�P��o����γ+򋭐E���������5�l�����[�}�4b�;�Z��!~�����~8B��Z�_���B̪L����Ӑ�p(��6`�C�.��\ʺ�v��R_�2��Yx_��9�V�/Gl�)˵����s���f����8|�ʢ�pz��8�_�nd<�V��?+��͢Yw�K������'�a�����=���x�sEDn ����s��Ej�_m;W=���/����^4UNC�f%����W�/û������?�m���ɐ%t@�[3}�&)�:ɗ#��eC��du����ƜQ��6����@t	Hв� $_M���p1�ҖvO|Y P56]~���ve�A_c�g!��5����-W�wH~��?��2�wL*��r��QCuh��3����0XliM�$���<��g�$�n�AqQڨiL��@$���#�R�&7֝�j����^L~V%��o%�)H��5rv.9�����mЅϊm�t��GMإb��h��6m�g�K����Ww#&9?ѐ����#��1+�I�3�>���M�8xzq�k71\��~�I�R��?t�O�b�j�l��V��8[ِٮxK�L�&K�C��uQ��,�A0/>$����c��/q����6R�p{��C�$�BZAg'�> >
������l"�܃���t8��UNi��$:p��DV1�@�|�E{�\p�j��m���A�^��=��DRI�(�7"�#����6\�'f��ܲ��+(M��>������ˇ��L��b߼�IC<=�T8[T���?�دl+�g��,�Id"�����p9B``=��/IUzE2`:Z��+�+�:xvG���"X�?�{x����B=���8ib.�K�0ί]�p��t1?��O]~|w��HYE�ӻʶ7�{�p2����{|����3{�5 �"AQ��1}@ ����5�]�>ߐ�I�{!���Z����"H���?���̖���j>�}����z��$O�8�e�jb ì�kͤ��O�mmh+g�������r��Mt�L�mtT�}�[lc�o�39�U��L�J#z-|MoaI/=�������c��?����zP���6eJڲ%�m��@˟SOH ��5���ѣ�?�
�zV%e��7�A?���JH&����&&�gyO�'00����)�7vkо�q���w��_6#M�uډy���{\q<�?�������@�J)��ob�͑'8��䘆��E ^dN�ڟ���HA�v��������Z/*t]q�*�ZQ�|��<\���GQ[�	���Q[=���4�O_�!��]�1@-�����gT�D;�=���梅���-��8��N.�3:��$_
o��n2o��ds�o��f�em�w(ߵ׌��
.f�ګԦ��-�]���-WE<�������>#r)盈����:(zAU?<��_�r�YV�����Ai�V$�H��ܵ��I����h>�P5��X�<�#��^A�S� ɑ!(�2�*r�׃�F���-^y{��gŰg��#j_�Z���B.�j@C�:�x��i`�;����H2��Ʌm����� ��2�.�fJDݯ��X}y-5w�&ع����1{a��!����J�h߼�K<�Q�r�J�(�����br�j��/`��l����я|��_om����~�찏�И�RAm"n�!al\�7-d���p�xq�cX��������Cd�*��V�K�"`e<(����D΢��חa�k�����q�<:���B4ɏ_��o��g�Y�s��$J,X�5�I9��72��^��1�.�I[�)��a@��őT[30N5�.���3�'�/���3�W��Ǧ��v0+��v\�mg�!��ꅼi�^rM%tT!r����А�?s��J�ݟ�Z������G(���������w��1�1(ؔ��#@�B���6`"Hb��}�ӦcL��oc3��ƪ�Q�]�	]�c1Ӿspip�7�BՈ���w��sF��p�7���v��!�_L���_#�謫B���c��#�<~�
�G�߭��nH���!)3"��̀!ְM��ͻ1�*%��-��.j��$IzZn'�d)�]�係Т2 ��4�&%aH�'6(��ll�驀4��uN2o���/L���F��}�k��IQ`xcm%n�?��%B��zI=� -`��r����i ������_�b���):¤d��K��G.)��'�ەg�d�	�t�O5BFن?0��b�,���;M��T~�f-Զ�y�#a'�V��3I�I��(�F��&��t��t�z9X�%��j���l�<yq��d�wMz(���7�AƋ���֩.�^4��nJХo[��&{G7�.��"��ӕ��Sq�dG|9X�f�|x9=�3)�>'�{�=���(0ړ�~���|�Q�I%��gpJw!e����5��������/je�.:@�-���0ezm�W:�K'���X!	Y^���+�43$�q��c=>Bg����p]��`D���A*��Ɩ���<��� �n˫ټ}h*\�@&���m�VEO�)�h�)#�p�.P�j��t.��*��[����*�o�z�ƽ��=�3W�4)�;_�p>��5�yD����u1�+L�饧&<N�oy�t��:)���oY��\C�^Q��g����N@J�M��8���>��t��#݈�T"�#u�."7��ϵ�)-劼������i��@び��@�tQ ���|�G����H�2yh-R�pR���u)L�̴
wFݽ�7����$	r��H#(����{�i�E�2,6 Y/;MmV���lY4*�{lj�l_��Yӕ|a*�owK��ǯ�L�|'�0�ځ�O��$��c��Pr�����6񪁮�x�����^��;����Vz��{a��z�?�Q�-�^j�8_{��-{�,��$:������`H�v���t��@���AS����+B�u�BK���ʞ�({yr#g��?B�&e:R��UI1�u�=�_��ˠ�Q���3�Cx�&1�&�����,p��/�i����}x�W��"A�����XHa�}dH�/CH�e�RU�묅�<�I�H^�DJ��Q��6��q�p�����{���gЂ3f���_. �`��3�\5xd��8����!�Q���2W>�g6K��Ј��M���/�@v�N�!��&Σ�@�)b�eZ�B���qt^�3Fg�:�7Z	���(մ�J�:�nm%��2@n�%�q׿������W7�t�~�Qd�R�K6~[f;@-�JO(�LS'�$�z����|g �����k(2�IR�	�fMf��ޯ�YHj������1'n��O'X|�6��'>7)�xޟ����UZx�&��峨Ꮇ=�-kTYE"�-��*l�C�Һ�k�=4��i^��u&k�y�-H��o�{��9B&YYQ/��G�2pו%')�egW��YBjR�T��� ��?�m�������h�:����^�^M�a]�K>{���C,��'U-ڍ���w]�����Ղ��6Km�����,Q,�e�]��pgaIÇC�2��AQ�W��(�b�sf�����۴���u&�@��3s�c-�/�>��	r�M`�x{~[�7~C5�Վ�K��e�UYi��PF[7)��$
�qa�^��(����B�����L&�_�V�0박@�\��p���X�-}h��(�xE0�����m05��=56#���k|赋��^Ǌ�vb��{<�P�oA�\�Jƃ���������Ø�y��H'jdO7���-�i�PO��͠�M��*pb��b��0Z�G�/ͭ�r�~�Z�fZ;�#'�G�~<�X�*t�7�$�r��ap5�UR�r08Az]�{� ������u��4����[p脦�a���Pk�d!Q�|�L�|(ԔAXCj5��ܫ�K�����NX�W�(g��s�C��xH��;*�5�c���q6Z}7r��/��z=�=����)(e:�Y�bԑ�
s�̺���e>Q�*�q��=�s����bp�	�v!�W�=����>{�.q?i��������%�
&V�S`蹪��s�6Xo7����2�%�i�+9�ΙT�<�9c����(^��	��R�[m��$S�9�m��_J��5ׅ��~�."
d��gW�F{B���6t>�X�0`����^<A�GӾ�N���T��B	᪂N���� [J��q���n�E�y�H�3����L�Y��F��̮Cx~N¹};jtY^�d�#��Z2p���;i�X<,�?�s��O��_0��Y}0��Ͳ�u���5�n�2��&�1$t�y9sq��P���" tbV�Q�\	�������k�����^����ӯy�v[.%p�2�i@BQ��:|���û��3+��f�}l������\�vgF�L����V��ʒ�aМj�J^ֶW:�����D�{��B���h�讉�B�l(���*��+��#�Q��8c�S4�R���]X��v@?�'_�@�׻�K9�w����[1`sIP:8�I8���9�����	�P˫!��&���L6�r�%a�}���E�@�-m$l��#!� |�$��hQQ�ݧ�
����lA> K���)�{S�\N��� >O�����/6���wi3����S2�)3CP�2��g	��g��
+�eR�i�蓢��$Ϊ���ӋbJ��د����x�1NDu�.W����ޏ�,���,��G������G��¡��`~�,x��tK����]<'��l������ȹ׻.
,Xvl�-� /E�$���s[���7no3�w�/�~���r�m��,��$���o'�ېV�{�ق���H!��(ӟϲ�֭KD[=��
���;�JA7Mir��g0O�t�l���a��k�.J1� �FY�&M�g��3&��n�Rf���h�H�Y�F�A
����Ã��l�C>�:u�6�5�Q�C#���53S�O-8H��[�@b�Kd�Z�C��r*'l�G��e.����m�PXa1�b��e�b`�� �L}��m����#�x��pPi�,=�lj�7�>k	�|��	5��+d6J��na5�Nn!n�SHk�����^�3�O���'8���Ɠ�J�%�K�s�jdW����|R�ta�v�K��t��IO�Q���m�٥� ����(�p���j��������T��5�.��[�Yu�����,!�(�����wn��(k4�_T��#AC?saϋ��޻N[��#���m�L]��f�/a�ô�XQ�ik%��C8����1O�6����ۢ���*9�M��%�x�?>��sUǈ�'B��0���:�����KM����N���!�f�1�YI���ŋ�Q����0Ձ�;��c��7܁,19�9���y5
	���|�߿:9@z+㯩p�P��:o�Pu\��6�����wT��l�d���e�l��bz)VF@i7w��N��~�ȤҒ�&1ͦKŮ����sYa��)��(Ki>f>Y�����C;�r��R���4�JgB�5h�XTe���-m#$B)b}e��;���
yy�u�-��u9�I98lW�?�ĦI�Ď��I��$4-f���sSo�;曱�C��vC�H$/j�
�e���j��p�⒎Uˏ���|�6�A��Wz־mU��2{g�Y�՟�3�� ) 7g�l�u��%�C�
�p�3�*�����:��R�y�&,��dBy����溬pg�:��7�T�cs�9�xCe�X�?E�JQp��)0�ǆ���Uٰ�	.Ѫ��a_�ͷ�����Ҝ�₰�"j�/�Z�j��P�$�	��`��T�n3��y�r<dkN2�J�#�0�t��N�t$�!,�ZF#\V4z�#�5v:i�]A+��j��r˙�{��9�o�pB���;'@�[ �����\�-��4���ODb��=���uQf![5��]��%�xnt�	�< D��$ڦ�Q����_���7iF�dߞa��8��_�?p6m��7i�m]�3}�w���֩��u29�z�$-���/�x��!�dN�yWs?��SO&�ş^��Wq�/��x���|�B�f��X}�}SA�@o�۾��?}�ټ�Lju�c�m�a`_1`����>��K��� �Z�}�@ސȆ�¼ �m�+�	�N?����� V��UBnVq�wK�������ɨQ�7e.�B�����6�]�l)��yH��˅���xJ@X��r�t�<����Ý�B��ɟ�ֺ����I�Pig4�d��A��lqs���~�4q�Lk��a�꩷K�!��#Og���Ӏf�a�Χ^{�7p4Gd���
beܡ����I۶�4�tx�G��a�!��r��LM������[���⽤�p�
h�k���M�?��&���`�t콂ݍ,��7{��i�SExa�%�z�A�)|�RH���%��aR�=x&z����}�h1�l�^�?��H{��0�����e�MJv����o��3��QH�b�C�J�#�c�3��_��$�:,���:���l��e���U��t���Hy�E^��#�z<^-3M"����0<n蔇T>k�A�lᔎzWjѽ(���}����D~NqXϔ�s��:e������M��T�ۄ���0>-u�����M�$s���c��qu@��DPB�ޢ��
�( ����=� ����#��u�	�dsmGD��Nt)fZ���Y�<���L;��=ޘ�IV��'�edZ��5�?�ba���@�NG��/������z��f�U��M"�Us�oy?�`�$h��Ѫv�����"�$Q����{`ŷO9��������,O�d�]Cg�y�/�<g�/��L*|}q��(�%�Aj��Q-�7�����w0�ǻ��v�d?H�с�W���L FȕC��.�'e���F$cV�R���D�5LFn�Z����熝f�[DP�&]��;���>�&�L/� ӛ�U$��xΚXʶ(@�Z�K�����ܝ�8���<*�7'�-����_>�0���n�E�<�䴢�z�tWK�.��`�m��8����H�nS��>K��N��������cc۴�O9s[��Љ�QD,!��޳�hA ���%�gA%�S�w�i�Pp�9���6#����9)�X�0��!�zwb�	��Ǐ�WN��)s1���|^h���8X���<?b\9"���n!'s��2�������NeG��X��j��B��x�oQ��s��_����Te��hT�X���3��9���D!�u��e���	�������%"
M�c�IW�dr�%X�g������Ihߗ�%�� ��7N����O��,Z_�@TMR��޷|�,�GbOh4Yx]hC��vySzH6��i�ؒ�w: @��y�*�ӈ���,2œQY��ga�,��vQ���.�392�#}BB��-^V���I� <�Ps�`��q*��Ȑ�4�]YK�^����?�~{4�Z��\US���hf�����H�-�LbQ� ��"�g�ki�{���[go���p�o��A��xDZ1��Z�1����O#
M5���(��}��<�~��!~{��a�:��^	�>N-�i'W�b�-��<Y�y,�C��Ğv��N`l�EQ�1�|[v;��TẾ|�n[B.FkeOm\I�&��6�I��LE��+�0�p{⿇��`���#%��<��d:ET��^&�C�_d:k�X���:��֠
s�1�FB]�;��儽�f���_̥���m�O�oZ�ɼ�H@`?R򵵺M��:��������F�z|g���q��Gv��p����-�~��꼫��v#>0�u�>��w@>�����Iՠ~����c�'�=1f��
^��ʅ�}KZzD#H����'n��Q
���2ȚZ�XY�sm#���b��Ʃ_,�s7��:���h(^X�1J42R�����-<z��D}QtB6��|p~��$��ȌuD�0oߐrl�WnGg��3� Y����4�)x���|�����C�����@[�.�j��X�l~��C4ʗ��!]�P?�PfO������?��f,/0��F�N3�zf�]�4�'-�x�@��Yy;�}�)��x���\t��ى,�fˣX��wSM��,\6�]��r�b��{��k�@���й����'���J�娒�_�߳J&�Qu �F��/$���:=TQ�d���*�v��l}���;[}c(��h��hW�;��O�a����t�ܳZ�rBu�%@'�gw}[K�"����M
2y?h���BL�m����@O�u�a�qK�gF��v�V���4Rq�>�`�^!��L��{��.���n�/�x���~�s��VD՚Vq�9} �DΟ1�ʘ�G����ňW�)������	`P�����A����l1�^q�5!�j&��:Z(�w^R
���6P���s#�����n
��劓��!`��7��9@ A��R�2�峤Yz����o(���A�)�����ˡ.���SML�KaI"e2��=�e��F�)wr�4bQ:��&z��A����BE�T
4	��73='I��P��{�'����3U�|�����Ў�T���R y�(�o9���8粑7;U!%zy�,�Z�,���I�������7��E�-��������	�u���L����R0{�G��k�@����I��S�f��S�G�ǵwA\����m��<�wĒ��Fp^'�,�+<�j��h�u7��?�����ވH�a�J��B%Ե�f�m������O���ޣ
V�q���~�iQh��;����M�U�����h�m��=�/u�� Z��w���
���~�E�$���Q�4N�
<��2�ǂ�f��;wL��������D8�0��� x7+�w��E{ɖQ��vG,\�7��5��!�V��Z����3n2��K*%��@��6;z3(l��7\��W%�/�#z�q��b��z2�A���%��[�` �B�)Y���{�9��&�V�et!�@2�@ ��.��ī�c�`�w��rp�����!���TyP��[���,ҵ�sP{띢>P]s��^�G^�D_�|��0�N��Y�U�FǠ�ߖ�5'q+֍?#vݳ�ϡ.�Aq�����U^��W[Q؋H��П>|��Vo�p?��
;��Hg�({�d��\m!I��3��-��z^�Q�"
�
�SY��-��,�d�Ⱦ� ����{�5�n~���g�o����1}�)�	�+�鵤��N����Y�]����j�1RQ،X����t���rI�2me��0R�CԢ���ZX[��`̦�����$�JJ%�˗�!����R��x&�E����Z�AC`OY��Z�z54[��1��u*=��Ca��