XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���؏\�eD�z����A=���pe6D()vyj����}N��p�j�S%svY�We���|�[;�]嗲L�X `qf>���E��0��� �s�-/k�fy[6!�oܢ�)��uy��Y�7�#����q"��J��u��{hD������[���)c8;�E��K}A������͋e��zfw�a��ԇ0�I[H�)�`�����,WR��q�����kH��KF������-�����H�)��͜)���3�(�/p+NTtJ��o���q)�8ufo0hxߨ�Y�"�<xL ��<�\�u��D\���o�׾L��N�F�F��a.Y-,M����7�҉s�� Ta�xh:�� ,�����Yꮦ�p�pr�����P3��}�B���߄P�!�vt���./}�/  �Y}�(�<���۹��4�:��0�m~�QP��_�T��t�D�h�2�������?��[�Y��%�.6p�`R��"`��ʌ�cQ}�W��@J(��\ꞽ�y�O�k�Հ�S/��Q8��a]��]�[���j��$}�Ǽ���+�E�/	ЪOٔ_$�	ݔ��âFᨺ���'�ݷ��'��l�V[mB�\VZ8��ۙzF�]� �`#��j!W��X8$v�4"p�|X5�JP5_J�m;w-���4�k�,�cT� 0b<����<��/��¼]���ZY��U?
��ĕ��-��\�O9ς�\�.�
vskG�ja�j̼5׼��8�:A��y�x���'�XlxVHYEB    3b09     f80��9���~�/M�g��3����ɴa���\[�@��+�2� 2B2Z���w��lRT����(4��*&cd"O^oY���69-�y�yР�� ����N�����#*t@r��5=�M��k�����$@����,ǀZ)���+KG�9%�5��3��[�������1zC��|�E��댃:iF���q�[�YAY*׿��d�Ag���c>{DL#�l���3'ؽ���Y֯F
���q�ܳ���w�(.����k���`�O���H�0-��9@m9��d�|��cZ,���D�`I(m����CA���c �]&S�M�dc]��P��l^F����π�Aj�$$`6����*b�KG)2MѲL�;��|e��Np {LT�r¼u�h
���p���W�ӫܩ��μ1j#���g<Yґ�	K�����F͜D��?H%��v��B�xFWε!C�J�e����^��x?�����Bw��5�.E����g�PzI�W���C}�����}��g�y��6��J��Vh�"`	�v�s�[� }��D��9݄�*�]]J&�\4���$aH$�y�֍�X�E�yx}֎2`��3����6�����୬�	A�Lg��U�j��'�h��L�:�5.�I���� ���۔�~�9���g��'��9��#��X���w����zMQ�v:��-W���DU�m�Փc{T�?�ì_�<���Ӫ�kAʁ�5ی/����������>
ſ�܀{�6?�|j4���5�D¨-Z�t�T����S^���=��a��, ��ba�4���6�z�	u=��=3����>G�,gu%!��~��X�$&��?ITQ��wD�D���7m� f�[��D�ͼ���^�O����~FJ_�����N��ǃ�F-�����Q��l��<��fU�f�VBzUG���|U�D�c�x���־t���	�E�/�L�z�D���
��;���$Bj�ռ�� i�'̛���I^Ը�K���k��K�	�(�NBr��f��Z��B����N4����%���v6�Q��Q�4%8�~�!��f�уֱ��O
�HT��!�wD����8L��d�fY�nݤ1�k��%�tkn�$ׅ�v���'4�]����[d������p]Te��8@{�c���z,��C&�;5�9�U1�~]�/���w k0s�W��g�e޺	�Ӕ�a��.�n_���,�Zℸ�>'��tA�4C�
S%q).��؂�o���m��e���&mh*���p��6�k�زY��8%(uF|�6�6߽z���	��p��y!�_)����	��t�[tIy(���7�AFk�p��q?_z�s��B~f�$,ꈺ׷���K�~i�XJ�ˍ�
�^c@�C��T�Y
����Е����V^��m��K�5�TQV2�)���&�go=Oؚ��I�ܨ\���b��"�F ��a)���w��.�$-$�s��n�7�BF6<z��KMS�$�\e�J���^�ؠ9�
Ф/e�?�~�Y��x86�s��@y�U�V�
L���B1&ڌ�_�hj���/l�=�lX��/���Yu�屈h��*`��+c!��m=��S;NP-o�Nin�B����}��~5�.�q�H��G� 1-��&`��F�����2�d >�V,Xn�v���*������7��0`��O�u/�vh��Q�F�$��>�9�Fp�w�Wnv��YCZtz�'��.ѫ�;"��2�iի�rɪ�w
,t��Pv� �gz�:��%;p�Ϩ�ϭY��M?%����h���%^f5;RR�kA�����/��u��XՇ�'3e�y��+��O�:��I���Þs�HTY�Q��E}ݍ+�b�p�l��%$�j�����������Yg�t3�e�F)wwIt:�Q]���l���&��W��J�w`>�g���|H���Lɀ���Cn���@������H��hb��NO�,z7Gû�{�xA��پ��_���2��H�'�2�uN�1Mj�b�1Pwmg�֐HF��$soֆXOʗ2�����R�l��7_�ctiTJ7]��;��J��vt����$�j�5�Mhs�R����c�Aa�����uy#�K�s�MN�%m4Ȍ��,|#�3H,7�!"[����Q	�(OJj���H{�쬧2���s7��Q$"ଚ,��'�.����Ћ�Y7�r����y0 �MW�Hm���8��t�V��z)I�#���|\rH��֕��V�ܓ�7Љ|8��ˏT+��})-��@5���9��Ϟߒa�Z����[T�H|h`mp��7\�=�+�K�?�8Y܆�yΒ	Q�@8�ng�����UK���[�f���1�jv���j���$dl��Y���]E��6�}C1Vُj�Ni��&�>,�Ո�FH����;�3��k"s��B�ӴQ#�H���v��Y|��%�P{TN�.q7�T�Ql,�R	M1T�y�ꏾ�=n�|�vw~�@��i�r"�	�a���6DPM��}�0vz�=�d'���8d����&�
�]���2 ��ë����/��1(�ÃkY��X㊂�i������X�6�a���.���	l�d�����$U計&p���psZ�׋x�M�V�;v�E�_ՇV1|�%([��'�6�p�iI��qk� �s߆�������S�$�I.1v��]�0B/�d�M�[t&,xp�(Y3�3���T�p!�; $�\���.%��p���wj��d��?�J^�gӱ aF�� ;�	�0��L��<L�ds��P�so0���z�?N�����n&l1�[��{�iVԿ�7�̟�6���.�Ƈ�;^nm����YZ��f�)c2/bC��s���S"���HG8s��D&1��D�F� �}{���l��׆�D���`�	cuC�v�O���>Ю�z%���ys(XQ� �`��V�}��mԒ��Y�A�<.���X���}��q%��5�Y�!��'���6�:��S���A���U�)q��F��Oq��dE��FrJPɣue��ӑ�!}�t�Xy�b�D޳����'rR-���(� 3^;c� ��s���"�@� �릞Ri�a�F�-��E�Jm�X P�ɊsG@��^���բ��ע�2��,�Xo�*,Y�q�&����H���}1��^���"�D$���Ba��8����]�$�t$<��w�c��D�(��9�Y���Hy�~�fGE���U�U�޴��c>ʭy_� 	��"v�1��S9yF� �B@-�'�Y��fI�$�#��	�e�p�D��Ĺ�9K�Wx�Xĭ56$�(�qKadOvi�=�@����s�5Tw�6�ꃐv5 )��_6��a�UO C}^:c֥�!K£e$�z ޛ0�*�]6K�&L�U`��I�f	��u�=v��ʹ謘�/���ð��G��7��&��O��X�~�ĞW�IjH>���ع��4�-��g9����H־��C	⁙��N���I�b�����b`~r{K��^�MT����� �h�@����p�G] aS�l\�(�дx֞GڸD{���U�5���X\T�#f��6��Y���v�ƣ����۪�;��!�훐�uC��T9�t�wg�@m��/�s��)aq�/���a�Ive��n��Y��'�kp�1i���XvZ���WˠU�hh�1�}E�e�T�T�h4_܄�̖�R��y�H��K~ՙ�U�w-��Ҳ�VczqF�����X���y���|\쩙��ӈ����w�m��?l���&�5�n�N�D�E��K~�j#�\?;M+�w�Rj�\��f�j���2�ѫo��.i<F�C11u��u��vC���efg3�