XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �g£n�a�Y�<�������&�U�����K�E�������#Ӛ˓L��s@�D�:�L����q�`u�J��ҰI a������ߚ��:C�j>G�X�c�=��+Q���7��9JQ���>���jk@�ǽ䇅��]������p�O�@@����e##&al�&x ���3��4�9��:!]rp��Q�>ɵ��&ˣXR����9O�W��Z�}oxJ�6$$�s9��c2l� i�D�\�v�cy^����!�懯K�#1#����s�~��.�3`).�%�t�8��(d��5���0
%�k{aԪ�㲽\����0���o玩_���6>�C��A?�&���XJ�z��p�8&�$$��y��[���ˍ�{\��݌�q���ݶ1�i!y,S�E��|殰��ԉ�����ǃp�/VJ����ܦ��e�����A5%T�]��wQoq~���+�̯��T ��S��փw�ߩ �9]fUi^5���t����Y�?����e��
����:�����@(L,�B�g�욫vxr�Q�3�bMj�೓ZJ�݆�/�fZG"�&Vh�����|�!H*�����J�Z�]��������G-�Li�B_�Rz�uD&)R!9p��iRpT��-��?���.��q�B	q�D�]��{].�6�#v�Z�ėEx�od�on�&R�Ր9A$l���]�Mpa6�V�ýk�d��k9t�%�����I����#�ƽXlxVHYEB     f6d     6f0)���)F9"�R�.�ܲ��1S.���(��Ilvb�y��x���a	:�X}^,;h�P�������!���3&ʚMn�O���'+���L�C�y��BK��*��d��Cc5?�n�����GHt�q(���|��|-;X���I��M��6#�E�Qi=z�{}R	'�au�����ӟ��I�nB��N&JY?�hF�_t�s3H��\vQ��~�>
{���΍�20jՓ��t)a���yY�Fw�p��.�Iy*��S
S|�G{N�Y���"��ԃ�EՊ�k�tʹyp�a[z'�3��_~�Y�9�>R��{3O/H;��������6^O�LY��SU7��I$s��;�}�l�'M������B�ï����7�Q`��X\�{��{c:T�`�W\�C�>3�y ��եPs D`��̑-�~
z� .qJz>!����ܸ�f!\�:��C�0�P�h/|�]�a,�!�ﳒ�Em�P��ܛ�r��,_
���.6O�s�f��M��;�T����|w��2ZxY/©&�3����Rg^�_U~L���hv1�$�3}]�r�[�Lg��n$��UXI�k�*�)a�Y�vt�z<��<jE�nd���0�-��g��J�gYFʬ$&+���h�;S:�a)��Ć�u�r�{��A�{A�'?�f�Y.(���}ʰ`�iYOsϦC�� ���$Z�x�Ҝv@*$��iO��q7+:;*�c���\q��MoQ�
�6�/G���<��Ҟ�{��8��q�N��*P�\@I�:&o�bÔ�Uo�"�r[�����<�@y���c�\�)e\LAD<�`2���t�vD�X��K5��y.���F��+�mM�M�)�5� �&���r���!a5#��l�,����K�}2Qḱ��ӛZ!d��U6��x�66�d��7ܣBP��&8�x ݕ�s(q���a��V­���������%в�1��墻�i��%y�G]�U��4K(��Bg���5KhOv���S$� DK8�I���� 0?�w�Nρ�����+=*�7<��-�{3m�7�d �������@��ޔ6�h�Ѥm>� njO_�s��J:�t��a�a��._Os�_,�����XC�pi�Ǝ(صp�"o�� ����A��1�����Gc-;����6���EOs$!oSËM���ڊ �ݻe���Y%B}����9�!�����������4���M�ݕ�k6瀅\g&|Z��f��+��ݙ疋s�ϸ���p�\�:n��R<���@�-4�P4D�$�Rc�m6� �^�uñ��q럌����yO�'�;�t��4p��O��wx� �M��W��B��o�Cj������84i�b�����.$4��̲(��5��1�SU`�(��]��C૾�!�����Ѱ�����~��ќ�DFr*Q@�cM�z���G�)^�� #�H��}��ؼ���3��[/�B2����8lE9���t��@��ï;�;t����M[��8���E��>�+�	؅g�F6�l�!�c�Ů�١h�R	� �$�.��M�S�B~�bx����o�R�N��hڄ��}��D��P��-��B�5ֻ9j�\�΍t"�(/l��hK&x:E����Y�l��X!�W!��e��id���=0��'	�!�|�yc�u����#{׃����"��ڧ��T���9�M��M2"[ל.����Ů��u�Ln2������w ���