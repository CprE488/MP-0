XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z �oOB*<���:hE�Vb��-��->��9�b/��ȡjj�A�����N�ˑ[ÄZ�� `�����ٺ���p��N�W��1�ݙ����1����Yd:7h쯙>�cf�eI���:9�J��c魀p��F7���%�W�f
A�:��v#-�JT9"����|��i7O�e�����2|vL�6�zt9�Q�	��S�' 3f!�/�u�H�UC���k�פ��֘��?N7K�I�K�#o�����!jA�+�����"'������Z�K$hDk�b�L�n��lZ<\;��T���\���j�kʔ1��E�;�@b/�-rg��ͅ4G����T�9�0�Q���Q��n �`�άa�*Y?tM@�@u'1����h�+y�eh�1h��w��5u��ϥ>�ϋ�+��9��0&�9ƻ�5�z�(Z$	��<+��LJ������q�s���ko����Wٟ9��F�Q�0OJ�����[?!.�
��al��_��]�G�a*�|���a�������f����y*,����j;ʞ��1�C��d�fv�i���aw����m�䩱�e�Xd^�Izc�ǆY�SA6$+�=�z*җ�IK����{��H2ņ����h�p$4_�5 �KCF ��$,�g��$L:t�H9st�j�<^�_c����'o����,<7����t�媲�nL[n\�Ȥ;V���I\�yTp��� ,9E���������f\�[�{SE�XlxVHYEB    6014    1840�,�͊���\81�HyN����E2z�����G��v�Jt=�He���Dmh#��gM��� �:r���,���\R�7���n:�&�Z[a�7�l͊��Mμ�:~��c�r��W@�<�Y�ϊ��I��ɠt��S�ܐ仁e��%���~g�]2��DE��G�Wc1����7�·�������*4���K��-�UĊr�0Nh��̘�>�ӑm�ue��V+�	|�����V�1J����̞�_�{�P �nQ�rr�z<��|NZh߆&ƾ-�}��:�1+���㨷�xS(蹯c�\8�a�1�)�R�[k�Y��͛Ȅ�|w�C�����![��N�&C�R�:r!�dy4�f�d�d#�*������0{�y�,a2!��ޗ��8���T���������;0i��}"��p���Qj|�r�������%�x�~���E6�`��wRϥ���,�IM�����9Y]T��a�eH��n��I,���ۯ��<���e���������-J��Hx��?�Fӓ*���j/৾9<��xSe��G�h^3���p����?t�%3���?j��gC�n����R�m�%�3�	b��CK��n�z�-��T&����vR������FJ$P��J;����D�˕�c�#���tş�ԋ���۳+��le �K8�Ŋ��|�Lpy�L���e��t��:K��Y� ț~�m���C451*MQjq=�E\�Q���j��V�lx���!-NӲF�'p������:b<��CnA�}>)��qi�@S2�����+D�G_�@��	��?)��j͡�IH����5�_X&/�BF[L�\�.q�U���R�q��4i���4fMR����(i�6~�M8�x��� Z0:G�-�Km�Kվ��`2;��E�� ��T�#��7r�}5Ο�{���q�7��W������^g�Wt<���{,p�v�6Q�z� U~�d��=��L�g�ަ��mg�P��T��Dڼ�Giˉ�&P��d\10��-�L��
���Q���;��O���Cc�G���R��b�����^�"2���K��R[� ��Q��U�,����Lˢ�*֏:{�^&b��.�Mм�|t'v��!ѩ��7�!AE�:^�h��|��
oK1��)������'+���%�a�^l!�
0��f�2�����6@�ǜxC����"^�������9�r�,�@0���dW� ��e�Y��z�
EZ�>Ӽ��}lbm��7�Z�:�ϸ=Ǿh�l)o���g�F��	��1'U�=��6bwm��azV����|/)����e�����k��Z��	�K��:t�:�L�P�"Ø��o��ņ�h=,�*9�O��qG3Y�9\��eh�j��2�N §n�m��u�\\.��	r�{����{�֬z��1���P^E�xU3�u#�;�6~@Y��=��f��v<� طpau�8�E��9HH��#��ޣڣ�'��O*�r*�j�ym���ɭiX�˒kv�E�B>�n	L����,w�Kg>8XYFR2�?>������6ETM���k�Ot���|N��
W۾y�y#������b�rs�}v���Ū�Q�e�� J=��d P�
�<�N����X7g����؄B �0`}D@�����Lz��R}�Ee��#�9���ރ��u�<����/NMY���q�}�(:����@��R�p��`YQ��3G��d)7�D�v�>�XɂR�GX��7��Z&��||��zP�)
>�e����DWL�0r�~WQ���u��vjM֎����w*ӗ+�T/0���͞�g���bje�>L��zƘ��uˉf���t�ػ�["󡹝�7+�~U�r>��c�~K����X���9X��"��7�X��t����{�R��9�� X�P�M��4��҅.�"�����{W^���8m��/	�b�t�$(ۧΛ�7���QeL}�m��.{�8�"Y	�G�����J�5�e�H��, ����������'�~."��r�����t�tаx��Mn�"�M��?�jo��#�^�7�����(���[dmz��ɖ�����^ԕ/��N+1��n5�E������.���Cm߹�pֱiӂ�"��:cQ�	8�C2U�]E�zm���N7���
ӷ\����;к�M�`�^�QwJ��~�߸���1�����6p^)-�K�xfȐ0C���"�|ۖA��f4��팉U�7��@��Y�TB������hz�\F@1UO3��P:i����Gag_&ؤ�K[q7I�1-���Ps �']�]�%(hʸ����:]����cD�kZ����7Q� �@脶D���@>�����(��9�m�*N�F����n�[!��4=�·X3*7�=�(i��10em@s���.�5��*�3�H����Z�X�VR�zv�նDհ���/	�h����<nW��b��8j�l~0���GA�.\F|��)� A�A��y�����Á@ ќh����UU���)n��4���nγ}�k�C���Z�uE�u{�����s���_1<ۧ��⃐&� N�+,ll>oy�+�`�S[ޅpQ�H�p��ʤZ�����D��-ԥ��Xƞ���f�!i�k�Q���:���p�%��#���o�k��Wf_�D닚�U�ꐯ�P�����s-1�S��Q�酞F��%K�Ɉ簢v���{
��>�]i�k#�c��+9���n�pVeZ9�k�ę�AM��/ k����J��9�zu�c�w���#˨N�~V��ܤ(�d�꘷�'�#���Wa;鴷��.�<�p,e����!�X�ʖ&��p�,�1^�}���q>䰠BE�&o��/P/V�Ypn{/�5�<�Ӹm� �r8�f��	��<��Wږ.`�>R��{g����t_|���������(uL����#�x�uGfb���@�������%��y�[�:��}��%�����M���B/�F�9\��h���M�Y���z��H�b�3���4�~]vl�)~���s�,��P�iv� H�O˫��'VkO�}��'`h�{!�����%�b�;|���	e�?$���n��u�����Y�eZжݰ�2`1�j<.9��3�/&��58�0�\&b9��pOx����?��c`s���Y�Cȗ�<�!���:9����;N�����7�,]�R�t�(��~7[���(�JN�m�㑍���+�ZFw_%Uf���ߤ(/���e��qxZn�F7��=�ݖ/�dDV����'� 
ojd)��W�mԼ�p��d�Y�q�GH��*���ڵJ�$ԟl#�I�7qS�H����0����RX���N� �k��scg�,��o����%���|�I98�[(M�@KQ�
�5�r�G�<}�@H�A1��P�{< û�E�\�3B��g_�����vH@����m?V\�S�mH�i�ZN�#���U�5L������t;���zPqs�n;�
�L���À2��*7�[O�M�N�����Y���>���J;CZ�j^�g�jl��j�e(s�'@�]n^4�,��%kczb�2����.R-���)w�����믚��J���HL��<���\\��6U�nL4���Z Hj\�����s���2-I?4�%�������l���V���"�d.K�;Ĵ��"<��I�z�ۆ�I�<��9OlU����[�p �]������|��F��Uy%�M�i�%S5`�w0)�}ڻ^2:9LiC��
��ئx{�̐Yi�R�-��=Ġh5�.@���D��9,�I`%��}>��h�kڪ�@�;��l�� �+���F�����H�[㰭߅�	$�Z�@�4=)F�YZ�����	VM)'��^���=a�䶒H�u���l�H]5�b��ꍺ���w'���-��Fց�VQA�[����t'+���rP�ٛӟ8p�p��j�Bc�����5PQU(�=�����Ay���Fxz���"%�u�U���R$\	��	�r��T�:�{���~B�~Te܌6�	��U�F����V(���_db�[ kA�����ۅ�<�m9���D)�]�	�?�Z�7h!�gK�#{�bx�����QO&�Xu,��:.uF2� �l�,nE�{U�>���G*iUh2�&�D���WAX�ij:@-��i3P�4p��	m�w'��\]�̀t�eQf�*j�o���k�Ά�
d-��z��]�ݍ�ҹ�A±��B��k�ƍ�*˘�pjhj��O��_���������4�Tj�^{�������H,C��BD-�/	��k��x����Y�FM�S����2(�P���o4�H�[#$�Q���z21|�'�ד��=�m:Ր��W7�û.���_�33ȩOqEnE��N3!�xAnb"x[��B�U*gt+`�S�_,�7[��󔆉��Ɣ3B�k3�h39����y&O#�c���u�N�?��ի[j�/�݊!m��X���x�Ҡs���̹�J6�;���&y%�MW�9�85�2�|�n���a�8�)&�t�/��%*�HÍ
ӤJp��n����I3�;�Y�@���3�i�	ep���G��
��,Uؐ�뿪(g���<�qFܝ�*ۦQd*���%>��;��,W]w���H�hW6?w�U����q�\&�\�.'��s����~f����J�PTj;n��� ���m������%�7��1[v����%�_Y;�Z-�d�l����RE%d(�7���#�����2@nC� w�!m��`㚇���({0��9Vī����Ll�q4�	a�h}դ�|O�љ��p暨7Zf��(�.��t��³F��G�-�7>��!M� s��N�h�/��=V儏{�D�� �8��]e�X[��(�/�/���/R�&��?�}L�|e�Ei�ȲuNUo��&��Uģ�C\����.7������o�������Ƴxu�l=�����6��>
',���_�w�����^�--5=e>r!�`��*�z����:����I.��8V���K�vpR�A�&G���z d�0>dQ�Z���M-�i���N���B^��ȈH=�2%o�5��@���{o�}�S�s:^P��K�����eF�u���W��g�[[Z�Hi�Ԫp`D͓�q.����(vL2[�3k���+x�
��J�e��r��|��aº�^�׭"�z�6�s� ��P���<hx�j�sҭ��!ѡֽ���x�|����E	���o�kZ�°�}p2�FX�yĥ72��q?�\�`�&��SVf��2 �k�0�>����Z C�;D�R��{���y��|���i��[S|B�r �9�8_����{�%d������0���Ϳ4��I7��)\���o���\[f͹QW`
o���L,Ȣ�o��Ц6F��hD�v|��3-E�t�GB�����v�'�A�!/H�ŝ��E�ؔ��
/�3�Ԣ����lY�4B6&��r��3L�(ܶ�56D�IE���S��#�H =���%{U�+S��;���]�`uF�)�&VG|R�u�Sb�IvL�x$�&iN�n�<z:��t0~�w�3�=��]�w���U�n��)<ߵ�I��%`��>Z}�Ɠ|���>)��v����߈ʬ4�I���M��M�1B�͔��l�����9��Emgbq�D����2�BU��Y)��Nf6>�T����C�'_\G.����$6��&ÎE�� ��:�"�4��}zOڒD��	�P��w�2��Ų��ɚ=,M��� p^����=��C��Z���x��z�\x�ǃ�,*�H��[n|�8^h� 4�=����N�C�>�$�z�S��P[�T��P���fR����H�ۧ�_�X��0|J���#���"�<�}�ߕ0�"<CHg��<���s�Dq&���?7U/�Z���˵ WCxYDg$���(�D�z��'#�c��:�|��4�4D$���\�	W �W��	�|�+gA�ŏ����tk%��gBY� 9i������7�h�ؓ�Bjb�P���.O?!��b5