XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����b4�`���8E[����@�@-H��'Y�����WJ��ǀ�Ӈ6 ��@��V7�r|�u�nV����z�#D){������`�A����ȿWh��뤧�|F��ҧ+Y�0��}{�@r�vSO����k��9��}=&e���v�X(԰�́2G�����Xڿ M|��n,�i8.C�u�S�C���C����5a>Tf��c3�0��;]��(.bYcG �5�8)�{O?w�_�v23��f/Z����O���g��rF�$�mܵ4������֚��������	Yk=��*�g��/�BD{�����ե��(�֢����s{׵n�-t���s������T���Q& �l��
U-�_���L��s"+��������@�}�@�u̧D�K;H=�͕�~�֍������9��`]
0���r�6�hv�saq_8_<ف'�ot{�������t}o�V�*���Q.gN:�+�apXC H����}��,cF��h5�ǣ�m���7����CkGA��=Y�P��Ĝ��ٯqM7;�F�pD��`�9���j���b�r��D_�=_��·�_��l�Ϫ$�@*�Y��In0%K��B��n-?X�+����V��[�n_^ʵQ�Z
�^���&���B��e��i�(��_�
�ۇ�V��eB���m�� bEJ
�J�@���^�o��:oUd#<�ʁ���2�]�T�>�?�F:=��� (���+�1z�S=6.�'H$AXlxVHYEB    1853     810�q��0�qjb���>�*��c&]'�g�/X�i9ZG)��Y3���8��^�MKUI.���1,�E%���	U(O鹈��.�˞�f�{*,�
rw�T!H���<�+�^p�IV�C8�y�p��ο0�aYk�����ah�YH�B�3���Kϡ���(94�6Z�f"�Vv�t^��ݿ�Wn1l�Ň��2& $8:�p���'h�!��>��%m�ɸ�8��I8����F�is�L^���2u��Ӊ��7R �/�3�NwCG�0<x��!F~\w�hb����}�i���!�"A��<я�K��XC�0�+�v��?���?��`��'C}��6P䧑I��C�Bq�Fu�r,��c����t�w����Rr�s���I ��hXQ\��<I���5��%�"��8#TI"���v��FNd��ee]m�i׍�t�����5�V�q�h�Z}��+l���|��w쪓�P?9�� 8�����k�	J�d�\�����$�V,Vk�u��U\��?M>��7_�W����9gc��4���u�yb�H���%-U�0�������bq�n�UM�^�8خ��s�3�p�T�a�%���S�U#���"ߋ7�H:��4[a�L��&�ŕg q�5A��$C}�ۨz�4BGK�d[ق���qs���V����6P���OYk���_&6N���e��f�]S�S���ޫF	�8����d_��� ���W��j�Y���
�
;��n|s*-P�VJ�zf�Zݺ!�6/�U5��4��U����|�r!��^dv���0�ʧ/G5�-�Ew<��12�`9�Wy9!��'���_V����n��]���l�߷hJ8+0eĖ�u�0G
����=�\�?�����XN��)~�e�O	d�paC`��t��0SD%�9r��w�'�s�+���������N>�Q��@�b-1��c/�J�1�w�4�ߧ��N,� @��1
��u5a7&���~�ȋwr���+��Dm_��;^�g�����'͹E,�9I1;O�{����^.�A�Tp�E5Θu���	%L甦Y��M��2m
=C&Wo��=�F����z�j��<ڍ{�:%4�{�C��.3;ʌ쒐Af���������!�K��4���扷�A�(|���U�I��t��.�Lt����,K�:�V�L�(�ٿg77�;~��0���"G�^Qb��?��q$A��nzXVQx�@ܫ],�ڍ�܊�/y���q���U�����SC�3��۵4J2CfŽ��.�M����KKx�j��n,Zq�ye�{��t�y��p�����O�Vr�Q��Z�m�(x�Vr��Fz��okf?��@/-V�E
l��b�NE�Ȋ2͏��R��)y�Y����(%�Q��#RC@�A� s;���}kB�5���g�����v%�f`��� ��#c�	� �q��	4B')����tTb�hN+۠ȡ���d�\jD��+e��R&�l�|ܴo�5����@�7��!�r���6͑ۈF
�>�:������]���QṠ���\��;z�>C���q�z�I�)-G���ݟ��H�s�S�YkG����@�EJ��}v`M�͝t��{��O�7Q���L^zc�f�ֶ{�L\��)sA����ThF{E�������� G2�U�HKSjd����������wՒ����/�c��P�m:]�⬍�p� ؈s�T����C�*ʬ��!�X�����r���w��]H�Z�=z�z-���>U�&uxC��O�X�jwgDu��J
�T>@R�J���F���Yn�t�0@-y��"�m�qLe�A�WE�{���ryJ��b���4|ۂ��2�dA���C��0%P3�v׼��~���F���K(n"��Mc*C�*k������R�����'����5 <,A�8���N��탌�h9���G�<��־t�w�-l5ۻ�ɬ��s�[�C;�u�vO��٢@m���!�5u��K�hz �57m�w�A=�@��Սm�h������,�,��