XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w����IK��V���[�#C���ϰ)lUk'��:&�a�����8�����N
�1"�Uw���h���� !���\�5���P
����T�;04#��M �al�<{��AF�����n����ԑ�Lo��~^B���}��~oTVc7�w�� �x���+d䳣+ޢAe��dǆ��ԕ���ȹ�|1|w�8+���D�Cl6��=�V��P�%ۂ���2�5,7.�v�8mt	�I:���Α�p��U�
�ɝ��X���ҽ6AI�8��<�$�a�T/#V���%ے�͆�60��l���X�d�%N�91�:qM�`P<����?r���{� قè������͐"���{ K���f��3�I�q}5B��\����T�s�a��/��RNr�����s��x�b�1�"5���Ď�W���f�5�Y��H:8��� �g��"
j�D`cg�Ap��fi>$]dI>�{ɖ�����T�`�����'P ʕ�o�Ѝ�c5n�?���{Qֵ}���>�+-�&�)Iv*���e�Y�cYX=���	l�1��K��ɛ�͘��@���L�3���sB|"���TE�$�g<�ד=��:2`�LR�{6e�
����+�`�������{�!dS q�\9`�f@5B.�ä�w��\-�k]P�� ߝX�4&w	䎊�'r�91<P��wo��B����H�j�u�^��E\.�=�Xl��LJ�}u|aay�ZH.|���F-�؝��삛XlxVHYEB    3b09     f80��J��G��������$H�`3�o"����d��+$��paay�L�� i��t���l=E�_v'WA�v�z=�vO���C���?�=�����Γ�'���f���ݙβ� ��*�����4���PR�E�� o�����ޕ̅�m����J�#�?���-���&T��Oٝ�.�~h�d��)���|}���9�J�ߤ�U?�Q/�t����$Ц�������$�ч�6���|/y݇����"'�O��Z:+(!�\�_���rx���&���g!�3	1���U�*��㪼:�l���d*�%a=���c7%��@T����e���%ۄS�.͈�0�ZǇZ����jmr�����y��e7��,<��ޝ�A#ӝ�����ݹ�)e���; 	aŒ���68���ʿ-Cv�	�)J�0̕@�v�ø�9i`l�7  /�:�ZG+��t����a�lL�{>�.y�ZA�B<��g�[pB�����DM�yL���N�x�$H��Nx��}�+�k��]Q���i����rn<���,{�����BH3�p��b��ͪu)ȩQUl�睊^7UE]���N���[�:M��vK��3dQ���'���Ht䵅|�n�3�5�t��:�j?$��G���XL�(TUY>-�."6.�h�fv���%�D��||�/&��<�;
�BX�I؞Z�9�a�}M"lF1�PmwU*��Qp,ڃ�'ƽ�q�z-n$��%<	�Կmf� ��j�n����4��[l#��@�L�g�F6F\C&K$��>��D�f��&����y�4�%�������z
d �O)-�׹��?zt�.����)�L�	E��J��_�M?G�����N�(�\3F D�H�p8[���@yW�d����;3�eb�G�����G�!�Xx����S�|�����G��"ּ�ifx���is�ѻ0� ����?4����tud���g2���^��* �~U@.Q�<�-�ɾ��A:Z�훌�#Pe�T�%4�|��Ce���,���E�'mQ1�%�C�j����/��13^�.���	`�+��\�FM~�<�r!�B�V%��[Wv��t��pĆ�z��{о�d:J����W0������Z���6�q�ض���f�q��� 9�]Z`������,1��xxU�R���>/�Wp����h��$�˹�A� u	�g�S�;�3�"��*o�:�ψd���W�kǺ�Dc%:de���C�1ds��G�JxA�<�j�bN~vMd��v���V@��^������0=�:���4��Qҧ����ֵ�K�uy�
��G2��x&�A�צ^/	F�[D�r(�����E�*(���qeN��kp��7���i)�g篥�m�|=�(����dm�ZN�V��E��:�˒�Y�}ozN�:�q�hW����ؓ�Cp�����Pt��04�0�̛D�@J3[!w����|pU��?��_s���$Δe��z��'`ݒ��������~?����Y�\
��:`�2�y�~"J��3��D��#Kpq��&v�B�̃�Sץq]�H&T��|\*��,��k������������A�u�E�&���)A�`yS�J0��l�V葴�-�Й���)�v��>\��o|�$���O�����]Fk������@��c�JS�=��~�>ᇵ2�H�8�d��"�g����}��?�}��"�"�%Ġ"��s�-�|I���U=A���n������sjP��WO�ѥ���Ķ�zn��1��6BF���#gr�]09:8�`iv���1�� �iE�T�J�'�œ4	���v�*ط[M��M8��*�	 Y���8�w��.8�B��B��w��JUd(�2���DJ��X���Z.��d�f_�cA��2��O��q �>b�`R��Kd� rڐ�����(�v�,ty��L�e�z�i��į�t��}q������%D��H&��N��G
3���é,�%�$X;� oX�j��3����@Aj�1�,�?��� ,�Cbicj�۸1s��G�F'�h�Z%@I�|�y e��\��9���.N��0���@b,�º�+�]	Vw1m����-5����ٓ��iPC}şP�f-R:o�hU�HAE���oN
we��Xh�#�K����>�q���y���5��"��~�d)�H�.6Uɜ�Z#6/�I� $��&0J�n��yՌ?��~�,�I��r|�� U���1���n��>�B�XEX���Je_@O��c�Fs� l �@��l��[��x�����6�ک2����ql�{��Uy�M��Ol��նaѣ��}��2�)�(��uy5@�R7\�)\���mjSu�c����&ۺG,�xo�u��Q &��U�Q��\��J�N�M��,*4�Er�ʴ�,Ւ��>�޶n:I�/ޥ���d��& �z>,��MW�UJ!0�Yy�U814f_[E�mr�>x��kb|S�aO�C��^���o �;���-.Io�_'*��_�?��LoF�MGWD^�2�jN��$u�ׄ��q����p�]L1o� �m���f�9�/`��s��\`H��xF�d{����]��4��1�&��<��X��]:�2�GI��ͪ��t�^MOK���U�_G�pͮ�>�*�b )=���mh�ôN������D2
'S�0�#�*Y���y�E0��9p.�P��� �7H��7��l��0�=a��/IW@�Ɠ��H�b0�]sA�!�wo��d����U{�4�4���Z0�w}�sVG�8�1�]���E������0F���/x
%�E��'���7�����z�����'��t\�(j
_�Y�h���R�Δ�='���n-p�ʎm�u��O	������>#n����m�Tg�������:Z��؅wqϙ�9,f>=�֜���f����ͧ���<�ү��
ș4�7|D��8����#%γt�)�Kp��p�>�Z󔓞�x�`s�Ӗ9�<혦��˩�� �9ؕ�;��!�ޢS]��^-���{!�ǔ��j,�0��<�����Z���)}��fk�VP�$
�3�'��%}��׉Q*��	��2owRf�:�R������Mz���J��ǯ��H,ܵ|1wBɐa_W�a���Q��޾F�[����oǉ4��U�!7���s�c�t�eG�m9�P���ȳ�px}�ڈ���6i\`_@�N�3�i�[������"��`O[�
*�P�߸�/�٠��W�F�l�3dX����*��F��n���9�;#b4S��^��{�&9h�u�����qI0;�,_:���9�o[�1�����8R8u����<�o���8�p>9d�Ll�a� ��l�.7y2�!���sasX�.s�Þ`�0+wr�[<%_����j��W,���J�=ʷ[6��	���~��g@�J�������l�}�%�%����?҂}��#�U 8�M��7��&u�	����L��E��֛��{o+��2����ή�e�0�����M���,�����J���D�}�~	�&�@IAمŏ��!�f�\��g�k�-v�Wѹr{��@�+kf�6��諝R�{�j�$����ڧ#�O�(�;1���]+��P���DOQ��� �������b�Z=a?v_�\�F%�O��V_�W�w��g�b[ƠT8���D��G�A*�])�N	��A,��]�g&��-[&����4�AoLw����.��hD�n�Q�!�!Zl���u7��TKzͼ�/�F�� ���ʋ�Ia�=�	�%�(��s0�?�I�|�=f%b&��l����4�o����)�:0^�Y��fS��[��'�2[�h�k��0�uN��/��-$9�;-龀���[I]�t��p