XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���5�F�`?�uO*�Q|��G�t�˛�eM��
�V�%GQ�"�Ȣ�N���7W��c&���� �&�9�I�� �HX��P0��~t�?�~f�_��DJs�>�Xw8��0lK�~���>Z5�#Rv��7X�{��l��N�Yy9�"�J��1C�ҧn��aن5�cf�(��� �U���=���=UM�ZF��{?����j�������7��8��
{)upݵI�t����P��^�hvY��C6;����A{��>cTZ$��o-o�O��h��&M���y��/����j �&��:�ʡ<X�<��F�6P�̾����X����Y����n�> ��ٍ�	��^�X���x|��\4���"�<#O���Dgq��R_Ԁ0�jw$���O F��@��>��o��w��xƊ������t�߾�ډ�����Ѭ�l�(��6@+��I�tP��|Ac�[�+L6fD�5���F��Ė	H�>D�@%SG���:�y����S��\�e�iRB�[H�w��ŉ��a!�dA���>�rv	�&���/Qr�[j�Ԟ��ڌ?����O����Qc�^c\�=�w5ŰX�>��:�cE+u�9�$,�	ے\T�S� �+�����;0	�����J���r����䀂�Xt�|4��"YV�����ؖڰ�.��!k�Z��h=���L��A^�;��s�s�Z�UV9p.��dU'�#��E�!�_祳�u�`�7�Ֆ���P�o��oI-�7o#�8���[�G�E�XlxVHYEB    3b09     f80r+��O`��s�6{���)�UԱ8Vr��Th5z�����7�+U>6#]�����$0��~S�H,�~f蠻!���>7�aF��I�H21���y�riݽ�C��v��!�#�67A�Y�ǻ25Mu���������(�ǩ��4������s���bQx�*屳�>{�HØ�u����Xu��c���_��G�5�$�uBL������V�X>��*f:����jM7�Dͳ��������S�x�?����>�r%���D*�hl5�/��2�5~�ɮ'�<���n9�>��S: ����W�6������2Qca�V���Nۘ^S�!��y�!Y�����.փL�'(���H;�G�H����)jYp9�ϻ���u�`��a1��r�F�#��8�׎�'��B�b�X���C��&g��˘m�&�UX��xұZT�����Y9����&�:鮮�MR�붧�;����%`v�.c�2���ɸY�A��VB��=�bV�f��
�_�5qnN���d�=τ>�c�~��7��4<��U�Z�>K��+ fEF=�1�g��Kښ�{�Qii�a��y�)������!�{���=�h��xY_�k�ߔX�r{O��@��U᭕f�L�(��4�Pf�~�O��H���ᶛ�HS=���I�}n�6Z9�mYŪ��E�׀�X������i�����ڍ%�*��N.v_�����&c�D�EG�v�����Jʲ$u��=[$�!]�� ��;��W�EdUk���Z���������#k�qBV�E~�H��2�K�+/a	J�Q����OD���ԓ:��0���� �y!���@R�E���^�A�^����s�Z׽�|bD(�I3��u���&c�GT�2�>��@V>�"�hTOu/٬$r+P7�z���ƙ�څk�g����[E���k��g��)n"�rqk���y�0��5����s�b|]3R	�%��D�]�%�����m���%U�mϽhL�rѧU�8w�o���l�����G�[�&'<������,PHI��Z����Uaw�
#��t��
4�ɽ$�ٲ�!��X��9
�o�ԝ��i"iLt�zX�=���(�S���`���ǅ�3\����b��p5���֟�̆�SN����J���~v�}�0�q�X"��n�2jv3ڡ��T�y�U�^�A�[�#v
L/��d&c���3�%�l
�M����S���<k�&ʏ�$P������X���V��[�����^s��v[�C� ��:U�~9��_��}"�Z�Xe� ŀD��} 
������߱OfK��Z+w�accF��f��O��f�����܅..i�0�� ?R��Iu�v;t*{>�z��X�h<Ȗ�tr]xNshVQ���&⫎�� ��Q<�_��^K��Q>s�M�Գ�y�N�^�9[<��MWF�������t���̭��_���P�H�E������A#+a��;�͇# ��1�d�v�'��*�S��MP��]�� 2_h�����/���j�_ g�nf9��H���uN� ��+v�rA��̣����oi�����2Fv���s�ղy��w��2б����|�߼	��-6��ж-���{��-}���a��V&���:�SzZ���;eU��:���ӛ�p�����m`���Rܝ�}������ɏp��o���Z�CW�Ͽ����&M��|�[�sۭ�wM��#��&h�y��m���c� ֥-ﲉ��>t�p���;
K'��W7l�/M.���w�0�r�A��UjߕR]�)Q*U�I�ؘn�5����B�2NzY]�`	��c����d%���S ��a�7u������m��>v��7�*|��h�7��͞�@h����w�O"X�|��,}4kq\�c�=¡7'��~�^L��,q2WS�6n�%-$;�����ʬ;�i<hil�j8��;���}���t��唨=P��uU%�
�����
{���A��qϺ`��+�DY��o�U܇HvT����]�셥?�]����P�4x�)��V�Uގ�[���k�׶���q��ŎB%�����1���K����3ѻp� D�-4����b[��R�z&��1�tR/)�ǹ�܂X�7sڽ�:�
]���{1��mA%5P�楗HA�f!�����	9(���[���6��vx�ro���R�ΊXVl�^�}��w]j�<ګ�`��%��@��F�5�M	0��ԣ�,A&R��.I-�R�4�x�r��*�?�2:�hIb,�6�&��}y��0�9��e?��vA���H���� �2�زHǬ?ʌ��lk<K}�u���Qe�B3�$H�x��HnGE|�`�w��͍%UV�����]G�[JRc�l���Rձ箤W���e��;õRӞ�j@��ʇ��m!3S��"%x�;��C����N1Y��Z�?�h����Ր`�`�M��.J��%{�\'r���;C,_����9;,�~]��S�]l)�7~	3���P8эY�P��̱�8Jp��E5S���H��X&��%E*:�;(��Y�(d�'���^�������^d-�w�O���R�@�3[�5������M��8Ƚ_�	
��������BIj=� �Ղ�$���;�\�!��P�J��(_S'=�Zt�
���)�b����l���ᾃ��<�k%���E�
i��� tW^b'�"�2��3bxmu�{x��)��S�Z�D]x�Tz����G	Y�!k�%�v|������P�ϴ_�w��B��ß�Z0�o^oW���bzB�,�;kDE�Pl��;W׮e4��#:r��L�.�cC�7��1O�Њ�{��;"'�2�Y �o��� �9ҩ����; �S��|��UT�1���o�1_	��I��`�����Elޭ�gT�ơ��B@=!�QS=��m��������:cj����"�K�Ia�z���L��ۥ@�ڀ�� ����E�3Y�L�"W��[-΢q0(�N�>�<zX|g܈~�����"�чIGUɋ�A�ҏh�b�ed~��24�6�B��~i���_/�!)�����F��,��$�ϲ;�#O!�J�� ꤓn�4\����$9���4�lk8�~�'���3��jw3���_�ϭ~�����kB�� �&�dy_>�l�4s����>�*��Y����v������\��`���ʍ7!b�qB&m�|ƍ�Z������dp^h�ʉ���p�
d��)٥{ݏ诧-SU���u� ��v�y>Vpx�a�	�4��\,��0�~�-?)���
�4u[�᳔ju9�T^0�����5d�EKɲ?N̳)L���[;�9�kwC�=��"��.I���s���gH�~�]�Iw�Lfbي�}� �9��p�"yG���ļ�^΄>2����i�
S���J'j}+*�Ϊ�W�G\yQf����	Tw�j��7�o���GX#��:�<&�[A��:1֛��",�g Ft�Y	�ܬz�DK\֖[3���$��m��M[��5���1�:�Ki���G�I��q�e��B���AYl�T��]�֫�6 �y�a�j_���ϰ�hl�����M�T)%�=�6��	^���?OX&v2�h[��r�S��B�Ʀ���,ewI�ӣ���e�[�;��d�k��`�o`�Y@���
zk\�:���e��y��J
�J�R�G0�p���%���V@#�=zZv�/��܃���r%4M���+ea$�t���՘�e�	Ӯ�TWf�ߌĆ������I\�#,��G�8��g7N�(z��_!T�֔W*�D�,�1��-��ڧ_�c̫��>r^�(��Md��m���>e^`jmx�*AIl
�x`�r�6�	��=��xJf�\m�