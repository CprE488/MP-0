XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����|Hd�s��� �:�\5|\nݛ��.?�Pj���w�[�"�PmP��R�vT�Ӟ�a�lyf~�M4��If�[�S@8�r1�`��
F,��U�3]{���wX����`#%^�i.@�Uǘ"w�%�����_}�Ů���5�|y�P��6������:�I>C��M�<>=�����^\ӫ�¾�	���z6Y?������uB|}�KwgQ�-!�|�{�X�O��5=K��㚳.��V��8�4�Y9x�vl����aNg���x��+���?�o�х2Pՙ�8#9>���uv���9*1jS��.^�UR^?3����Y^��s�u�q�`"�m���uB�KjQ��w��$9Fﭹ��&�.�1�q�[��=�<�%A�'2� 3؝�`�6Y�o���|�w�Z����+a�=���^�p1ߗw2_.\Ppy"f`�& yJHPM�c�*���:M �.���&<��f��%����:e�x逩��(xs�}�Tp'��ݪ&\_ofsVR;\�QFc�> 4#<x06u��b�D�ϧ����#�V��D�zG��/9w�����kN��&��L(]%�� ���zw���/��5x^2[E" �:��z[Zk}Mh�1�G%3���w�|COr
F%V�1w	49_̺�?VE�^A����M���"�=8�*���}�8#���W٘W��"���`��2�=!�j���qT"6�<�D�7�奷1O@������XlxVHYEB    3b09     f80Z;�ꏞo*LUw������l����)66R����2tl��^� �����!�-���Y�� SZ���EV�pm��!��6����M �!^[�8�4@:�>H�/�ۋ�U{�KI��r�i�G��Zc�d�h=;P���s��,��`R��z�ț��XH�&)�n
%D'�
�^��2�NT��d�1����K����$$�6��	Z�[;B���J�n�R�����e�ۇ|Ś��ᓲ��0�Qw���ըm-�lx�S�w1svj��lS���-ˉ�6�,�n9uR�W������̈�v�� 'ئ��J��Fb�8�7�:����oX�h��`r�Rc9��Sr�|�8 $�J��$]�<��T�@&��/{�
m�{I>�N68�o����s?G��=�l�N�C<�d<��=����J��_ ��q�Ǣ��V4��e!��-�[���|�:`O����"��-Cg��݇$��4���Nۿy�3wE�������	^�D$�]���0(�D�MBwo��f�~+3. b�H�W���{���3F�y'�ƪ2Jو/���~���R�?�q?�h4��6,u�#إlF�3F^�7	�?m��I^�u封z������Βk�i�tpQ_)�P'L[�ZJ������  ��Y�AC��$Ikތ�y�!D=�9Uؐ+��Ķ���}ܛp�P.8�\89U���~J�k�^�Àd9S`���%k�6/�����c*�8��T� ,?��� �.bs̠Ks�H��bU�c��ae�]m8W�<��V�8�>�EM���]�mP4���}�Ty�X\�H�t WQ`�e�D���P-��}n�s[O�\x�"qn�de��#���?�wd��Wȭ�t=� 	
h*��\��Xg���U�	���/�>cW4��h�V�[��.8˾m&�L�ڸZ�P!���� ��s�vmK�֨-^}�~Z�毸���I1�����S���&���｟�ڬ��hh�7�9�&Ȥ����|��v��TJ'�,yZ���D�O�66���hp���F(H���Cx�4z�,���kvv��y�q�V�mx�ט�_�'c�� l9���Uh��2�נ(�C�d�S���d)�����z*#�gW���i\PݖsW�إ7�я��Z�Ў�?��X$|��\&� V�| tH_�����,B�����7$��rG���E���"$�_����s�Ki��z8ty7�|!�{���bz	 ,� �	�Y���b���x�-��g�6�L���t2���v��2�#4��w���I8�8��O�yN� r���\��veHW�1�=�t����|�����z	�oe�c������ɞ�0fx���"�I�*=UwjF=�Y��(H�e��sP%���$;��u8{�I5��)o�0�����ۍt��VH�>݌(n�YU�&c���%ߠ)�"���XeT���ǩ���39�y���<�R(�G;!��?����+���D�Y�_�ʕ�᪎�^�}g���>0dɶ�R5?xf��I��B��ą�@�!�����~��d�S��������2հ����W�}���Pj��yx"�~��!�}�v�0Ct�F%^�k��W���me�sÇ�2%y3�'�0Dʻ1� ��r5&�s�&�@W���*ނ������Z�7���G1����{����9�ؒ����${��,ž_[m��"F@���a��}�z(��J_���ߤ2k��������>��U�~S�y�ӷ9%q�N���g�F��G���-a�țy0T<����ܛt�bQ;e�����0\��7��R3�%�}��uCJT�W-~�,��E\5G�:wcm80Y*��a,�y�`��n�1`�����B�w�R��������h.	��P<~���$��(`A{�F"�0�>�i�0l�A�\�77x+�@p3��k���&ޙZw���t���WJA#�Ѭ��K��M�����.��,�2���
k�hLٜ��.�K�G!�0&��VK;c��2վ6�Zf:lG2z k�L�L4�^�bP��T�������LM���S�>�zF�j�7e��X7Y6�j?<��
��r��ŧJ�)�OSX>� ?v�|�E�;���,J@�n�	����1?1�R��$.Fpqm��m�0m��9���6r�T��S���L]u-rutuR�B+����Ӥߖ��fJ�Fһ�S�J�A:,��~�xD.�v8���w{��b���~�zWS��
UE[�X��2e��(0�ĔϾ�a��}޹.���|1��Ar�������q�&�s��ʘ���D0�@���v���6U�tv��c�I��	氠S��D�+�M��f�F�.v��&��״������[U�=d��A��B,�=C�e@���� ��l<���n�E�_k�����O�:�x�ꁶ��2�žm�s��č��S&��:�ݾ��lእ��Y�y�4��H��N������?H�[���Ov���T��6�G&Ml�`g�摑�\ڦLs!��X�3�H��6I�g��֭�a��UA�F-�ps�EH-�{'�y�t۝q�uO��'��y)}���Y��rr�u������P�g ��M��!�?� ��SK|�����t�ʉV��$ķkM�ݙ���Ƹ��R͛9�:�x~>x��y�$T�~���_ť��|܎I��*���8L�Kl�|�LD�	pj��V�n���~�H��S��K���0�(��x'[���2ӹ���Fg�:�<.cǕ�c�����6�!� ��� ��?��ͨ�T��[X!��֟����%�0����HU$��_������論���_�8>o��y�9�x���](M�A�_�NǧkM$^�=��EY�<��F��߂.���?�g.�x��tJ�N�[��~�ǐ��_*��ئ!9���*	�=�}8(�<�8�����rCQ�����^J�>�q�hB-�v�Ғ�4}�z�����1�����%�e٭c�8��HY�V�U_x��ZA�x��e����9�g�cLX�Oq7�g��A�c3n�?��9�m7�v��G���p[�����&�2�4�w4i?ZRĈ�he��e\�4>��f��~�h�Z>�hs�ŭnhl]e|�h{=�9B���Fn�Yǝeދ���M����6���>�Bu���@��J�Ž ����,����y�|�^���7�����j�6V�`�]J�=#i5�p�|R����~6Hh�~�mVF�0j\�jɰ��x�����.�~�#&������W|?��Ɖ;�OSK�R�y�ܳ�v2h���[>Ɉ��.�<�ɴoU���bJM�-��t��iU���W)����G���E�>��V ����q���Kl�����yD0H�m�Y�Yth�f�G�	�/#՞���{An?8��`U�p�zxI
8�,�6<�m|]�G�A���wG�2����$�j�3G�#�si$�JRUU�* Duk֣"�I�#)�����<�
34�Sս��Jo>�vi�ή�Fh�`��9�"Kr�#H��dAv�A�QA\n����uF!�@~�z�FL&\9�<쫁`���}� ��\ ��u?yC�.N5G�I�����DK{�?��ԉ�����iQ�te��J�D���[!���T1ZQUNK*��8�Y�k*A�����N��_up�h�������S)����������ݞ�?���l�	�D��^�G�����K�ܑW�.ůs�o�.��Cz����Z���<��������$N�����තE]��-L�a{���ʽ�Y��p�@e�Y�V���E��y
���������@���lň�s�dg&g^Umu���+�����~d\@)[y��PZ2���DW��Y����!��/Q��Z�,ӗb��8 ea_