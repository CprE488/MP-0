XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���P�a���
z+�;��Q3�Yw�++�	B:<.�#Q�*l��1�$�p����1\nv��Gk8S���jQ\7̏s���sϛ6>�>���w�*vcwܜ�;��]$h�!��������bؠJG�pI(,��y�z�*g1^u#R�n�/�]�i@��&1KCp��J'1H�����G*ʯ~,Z�'2��O�>ܿ�Zփ�=�~=����k��I$��A�EU��eL�Q�������ko/����e�U�S�U����T������s���@�T�QX0��rUꖗ�AH��3���P�i��
�H��C	|��r��q�I��i��s^#!{܂q���z�[l�H���i�Zaq�ꧢ�Q�@�[M0-��1�Y��ci������΀��14X�I��d�a^���?b��� �`�@&]R�B
��ΡV��. �O@L���f��s�������2����G��&�ލ�z��(	"��lʹ_�!p��B��D������(/�pw 3��^.�w���┿n�����Ovە֍�4�gX�E-f+ρ��zF?l�PHd�[{�[E�&�6�8vZK >O@A>߲���h�n��ł�%*�+��xW���xb�ϕ\ص���&�c�{ē!��&rJxE=Wy���s��{2t)���nl�j�Ǆ�_3i^���w?BK�;F�AC��J��cL�׽,@��<ioU���Dd)���/[�^���� ����=A'�2��!0�����e�-ˡiXlxVHYEB    6346    1790j�"���Ŀz!���d�ܘ��`�}�Z�QH��ŵl˫����^	��b�NKu��A�(; j��S����q��?���V�WP͜��yl��:&!�^!�	;�~5>;muy�$YM�'c��`I<���2TcסRQ~n�OA8X�e]��!�����_?Z9bf�	u�eb<��׀�� m�,<�[��kd���Kʐ�5l�e�$�v.~d�1����	��G��*��}pT��'fS��J�g��H��e;﹡؎��!��
�b�ӹ$��{|��@$���ܖ4* ~��d���Cu��G�B����$]� �Bu'[�<��.?�4m���'#�:)�x���HߠE������a|�1�r_l _�!���׸�)�-�;�"���r%��z��O��Q}CӔ��FX�iD��;B��`7pg��o`����<P�^�^D�$L���PI�ȋ�a	��ʲ4�0aOִ{Sg��\Β0ߗ6�pRY�w����l��������\bu����f�*h(���W`����b��E��
��=�Ӂ�Z�2�ʂ^"�_�2cǲ6��J�r�V����cPq��F��}�����y/6w�<m�WE�WC�n30���KW�
9��\�^?<sH�z+�Y�k՚�KE N$���21*�@�:Kl#P2dt�3��Cf꠶���d��Ga�uy�Wc���v���|j�ƣ�D����<	�1MY~�Z�u�|ˁj����i3�p?�ަ@��$0/��Npm���t����y[�.�ה���
� %�R��9�Y7�s�f�$l�i�}�nG�i��"��T.`�C���>8�W��t��6��b��ߛR�(�=�G��Z��#��e:p���k�[�P�N;���2#Y��9�VK%�?�,Qϻ���
*H#�l��v�������t��&ȃKG����畎Ŗ��5���f��
	�qD��S�K(+qm�9D|��0�'ڏ�	 /���
��|��2R���-"��3c�_���H���)��/�vVS�EdOZ�H��3��U2���٦�;M/�Eύ� ��.�<D~q�6i�C�yѴUp�è��l��N��OT9gJ�ϙ�{�nҵ�(���B�3)���.Z��n��H�E�j<h�+����ꪌ^���av�������S��2g��'�I��v�)��,.��D���Zo����%C{?5����@����F�h �m�Ŭ
IR���
ҁ[�xh��+{�Dnyf�004��uV��o�@�yW�wǍa!�ȃ=2�6��6m�LJ�3���c�x$��L��ɛ3�_��SZ�:J!��<XEi>�n���t	�D=��b2B�a�y��3�´yo�5��=��B��w��G��=��������
O���G�c5��eu���N'<�~a��.a'��/sp���}����YaJv�5<^%�LB˷ƄB-�*� Hq'*O��3as��"��R�l��|p ��(��s�(Z�w�3�����HP�V(�L�a�X�o�>.F����y�q�F&�F`�o�!�ڳ�a)$/�^�m���ߨm���n��#��%7.tGN���jR(���b��1�&�n�9�d`�|�b������_���4.o�G����_�����b�l�25}d22���S7�0��*�Fvݠ_e ��hM�	��t��P��	�E^Z�ů���\�1�]I!�j������k'��q,���˼��~���|�U��Jm)q��!�(p�$�7У��?(������s��NV&�=���˸[;^���;8i���5��l��3f�Ӱ3�9	J�dt��LJ��Õ�	<�dq~TW�w��[���$�{�YYK�h}�����_:��ё��C�=%5��0��$�"�t _�,w��~�A٥3s�*-r1,wj�1z�h��O͙�#S]�o��r6u9�oSs�IW����� (Ņr��� l�2r�}�J��gQ�K��z�(hڙ��c����=p�˯+�Ml&l��K�F|&S�Zm r-�=B� ]9%?)!s�;�d��#v�y
8=�41���]�@����$O^�Mٲ*\޷h�9%��M�D�����)ʸaF��\�h$A�䃛T�-뇯�X+D�Ub[93���y�ɼ����u�fƖ0�jY����q��nc�,�SN)lO���d�A�\g�L��3�(�JW��cȌ�4Ұ��C���i 9���;&��q�a�O��_��F.��D�&(v�}�b2��ѓ�q�����|d��z|c�I�C��wN�)�ό�&�Oq��Q�|x�3���E_V����z��h�R{��u9��l�>\��n��_���St�{�j$:R@ӛ��2kWz�[�y8"ɣ?�5��l�v�뾩+��K�%=S���3�!^Ek����CQ@�꫃�q�!p��/*��<?��s }P�~�P��f�n�l����h�HZ�ۛ�Z�.>_��}XȌ��s�s����_�.L#8�G0������ _��uMt���w�V��=�¬�O)��·��Vsi��uR�~�e��m��%o�_�p��9�["�N��0��p�y3GM���^}���)ed��(���\�w*ݞ����|x�_�U\{C�Ɍ.=�䂕2��W����@�
b���M�`��R\fkJ�ڀ�i�Fhn���D���MϨ���~����'�ڢ��;���T�6�7Tw9� ��6��6o��
�B���gL퓅|5rV���s��m�SA6=
"3�_�k�8����m�a���.��� J�cu�$��g:3���B�BR�w�����8��[�.T U��3����F�i�o_g�56��v�0/�/Ά�APb�(�� ʌ�pS Ş�sL�.)����#��l)p<�N�Y�:��9� %-����<�h�#��f����^�k�1T^<�`E���;͑<���rQrE���I�h1��ZY�ݱ�/C8j�W-g��0�αaa��$�&��^��$�)��~�#^+:��n�
����ǌ��X|mc�<O
R��^�7T���.��=�_��-�OVU.7������.n� s5���D-Z��n@��q�QX���Ɓ�*#Ga�*тSu�(������+�.�����qy>(�������<EIG��}�[�R�)�]Fᠫ��"�8W$�!�5���-3u���mO\l^���%�ve�8�Pg��I�X)͠�KE�`��@�F��E�Vd�HsӖ��֨�q�E�y���&��+�fR�A��E��neǇL t̫�q�h]׮Zj�i�*]�m�}��Nc������K�6N;ȢZ^�X%�_���-g�1��O[��z��~n<�c(�ށll�	E�.%F���Cp��(B��¹S�vҸ4`O��#��f�aM"�N��å�UP�es:Wj��4�ir�ؠ��w!tʏx��j����q�m��m��ֹh��j�����w��z
�qz̹4����c�ym�&���d)?�`��-�af���,z���Ű�� O	�X�e�����mzrg��^���e����s<��G�4z��+���Y��6(� -�{��-��4I�s�0�ԡPk>|]�y:�Y��'��+L�ѽ.����q���$����(u��{�9��a�7G[�3���P�'Sm��iy�p��/W!}�YF)ǭ���cNF�K�nP&f���y^���4\��P�{�;�G��ìo'O��3�A���+��C�{��$�9�dEol�K}�^R��������Ϻ�����e�������mE��Əb�P~��$Ϡ1N�!C2�"��mz`ˬ�L���ۏ�;'�0�nI�cz�#NR�UL_�"�yA���ϕ���A��Ȅf�8~�=�D[z6�͂6bz������T�6��_{�9u$����	�0�$�/��Ź�Uv�v��S�vJ�'>�[�܃�d�l��/��{��z�[�G\��%o��0�ހq䉘P��W2r���0�ɛL8Ew{Kp�4-�M(Ta���f�7�d�_��KF�4�>h<sL��[��i�=�p�B!V<(�����DK
�A$}�]�;Xd�7�K1��d9[�^�D�^�MR��E��`�,ꬨ�{����>�0������`�#��%cΦ$Z_��b h	$��t�M��ZUs��XA�%翸�x?�iA���<wXx"&�鴮0��?h-o��� 8�#�Yy���6]Ȏ<_S�K͆�9�U����K��u҆m��L�p���2�Q,>��8~��8x�!�ai��u>�-#e����o�i����BG��q��y��$�3�voI˘1h:H��i���bbN�2���	i�8$`��#�S~��o�&@M~���9�Sx
��2%��^���Q���_^��!��������
����� �;���\��"!Ln�܉�,v�2�������ˤtۋ�"�x#?�QHϊ�s���G}�Fl'��wh����^ށ�s��f/���j|��"��0���)1��82�:�o؀�<�'�^b>�d����j ����	�3U�Aw�-l\Bp���N�g�I=`�/"�28���F�5�[|��@&�^�fȮ�>��t�F&�H����Ֆ~qʙ���!Y���O�P��>��?��=�$� 2�[��^��JI���2�Yx��~����,�!��{�pSp�r`vLP��G��t� `uڒv�ϱ���t�eg���'�M���cgk���d�ð�HY�Y�����0
>Z:�y\���J�����#�Gͣ����G{y%�䑟�Rk΅��~�ͺ�s>ȷ���3���1��@�ZLmJL���!��6��}y��R|Pu���e�j�B���c{�ݚ�����:!/f�,.dN��5����#.�:y*���)\!%8ߧ��<ީ�0���&��˔r��fx�ۃ���<U��p1�f����i������v!w��ˌ��^&�7���/G?��ɴ�8U��
�'��r��0��3<E����w�&�"�\*�������QĲ�? �6i��[�%�U|A5���twy;|��~��c]�D<��x -�0�$z��0�~08u���CF��Kf=�Ƨy�8id��D���Z�
��΂q�!}�O9Q�E9ل��*wq�ݳ��t��g�m7��E���[7 �w_zuD�sc��7X�`��Y�{� ���}������=�t�p9f_���z�G@�`a�Ve'�q6dSX_�+VU%ԟ^L���A��0f�)�sN�|���bD~��t���
G��3��'f�n�PP���,��|3Nn8~��Y����{Y�^{&0�u� �s��������?��-+�._���F˚��`��X���?��#�ׄ�d����1��.�\F�Cq6������'�b
�Kq|^RԄ�J�j4o|X�Op�fO�� (-�+������q�����dӫ���O d�˫)���$R�ɄhY�!FBL�5�PX��6��)nvyu���1ɏ��
G~��,�>�7���m)<Ǆa���z��C��H�!��*0���XE�_�b�U��HV��p��O�8�,����
�ɪ��y����P_.Qا�q��i�O�/�u�XBy��m��Z{��M���;��������JW}'��wGY�k<��37�L�!L�h�p�����q�g�Ji\s-��5���ڧ���!2W�& !�y�R/����[���smS��X=��T�c�����t���tg),>A�2��B�/��}�re(võ )��r�a�q*w�eE��1���%���(����Mw��"$M�a����v5|��-E�iO_aoyo�����l�����8�3p1!��$�7�
�]�(������bj!A_Ý�璖��~v��^
M��E�`^p�x:5��\���Ȍ1��X!\�+�n������a}