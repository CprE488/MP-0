XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��" /��Q���Y= �M��^h��?�.�H|�����п17�/N��i�8ׯ��>�x��,����o]ٔ�ԣ`�(�lզ�'+{4�ª}�������XL�K���	��2oϿG�(��-�["u����� �;=����Gw[�t� ���I�{�*��[-�m��&
����-��E*�i��,}
�f8>��;�t���;�s���7���~|q����ǛY��E�U�3��?�rq��'�C�םː��`s����"¥Y��Q�I��J�c;��K%��.�>w����&�[rOu�(E3�=�sL�e��aQ����	��K^ QXL��y��A:�[	$�AVn�0�o�Q#X�]�:l�>�P�@���6M��psUQ�`c�&�(b'�~�k!m�/n�ߪ�g���{N�Q�������c�˘WS�p3�[�+c���c�tԍ&�N[:D�R������z|��jb��Z��y��v���4_6Og�q˴[�rr�(a{p��������P�9�
�J���o�_n�5���8��W�ȁ*ь9&������,��h/�"F��6�?����zq���2&u� ��hS�
u��F���9���)�ö]P����G��E����-f�o��]�l��_����e��6�'d�E�pD�?�	�,�=�Z��:�:bT��v1���z���E6Q�
ˀ4 ����Zz�G��x` ~���z��\�),�J٭�����L�G��nS��R�}�h65�I�J�ĝ��XlxVHYEB    95d3    18d0���̉�.˃��4��:3�5�b[�d�ڃu�0�I؂�K����&�'	�HY�q�9��$�����w�(ЉI\�S&�N� &�����0��9���H�&3*���z:å3���G(��\ÙP����rp	<Q:qh^d�o�N٥p��$F��v)�e�׷_�P�f����&��
(I�,$��$�J��x=�b�w?L@�|�!a�Vy�%�� �
��\2�8�<h�9�0�	������|�d|�̻O4�u�������9)�Y@�C ��%eQц��p��v�&�7e.�o���^����V+��M���ʛ����[��]Bq@H���o��e!Oxv��̤�u�M��e'�����Џ����R���u؟�f��U_���eQ!*�Z6}~�CB��2��AJ��ڳ�/�<^��H'�Í �+���i�98���L��Hr�[�BO��ߘͩ��P>�e�1�]X0�������]	OB�T�&��-��]`rNl "��ʉkk�g�?v��㶸�c�_��]�`d��i�k�K�����gR��ze��5XG�0�.���X��Fת,b���Ô��X���Հ�.5��{����v����.�I��2�8W�e�������j�P�!J,��}b�qT�J�u�F,L{I�i��@�cq�a��Վ_g�gU*y���o|��K�@@%��#�F�f~9VP�=�f���^cZ4e�xٿ�;�b��)I�k�v'�~�����Z��LV8̡����d���}��ۛ�� ���1���W��eY'2�D��e4�SU�Z�<Ͳp U��,����$HI3��Ɵ���.6�	�mQ�Dm�A_�&D�ϳ��Ҙ.�-/8���e�~�}/��n��?��`�S�LaR5��8+~Ѷ������C���7c�[�FP����b��)�ܲL�B��9�U��LPҬ~��Ԁ��'t�j���|7B@��)� sG�^Q3�C��t�\\s��*i���Q���pNt%K��6��X��*����q,;���i��kp8��,W�&�CA����G�+�k��Z�-�%\��!�|�2Eb�c@W��%ى�K�x�}�]�>U�?0X؎\�o��� �8�v=ч'�?�II����GY_�~L�b�\q�w0'?�'~�4'	�ӗUl��J ?{���+4�� w�h���Fм��'#A6�*ęʲ�>�fŹ\͹U�B���-_��$	����7P�p�J��u���[ޝ��m�b�1��;ޱ�t�t�q�BM�5sYC�V�t�.���&}���H��e�?N���(zb�E��_��
����}|���B��6����~+v��V[f�m3\���|�-�W�/�����	��Y����9���4�"������?Q!E�"X�Ꜽ�AR�c�=��1oh6���]9��c�����ߦҥ�A������8���l1���@I&k{�����?G��Y����7�^���� �4kvU��V;�\x�L+�(�{�y�1�w�R�]F�*[@e oԥ����t�A�^�;V�lɾ��%oQ'ɚ���G
��w1�a_� ws6�]�؎u��v�yLq��56��;�v����]A��q����뎦��qE{$gY�/lt�$=s��3��a:dC1%��>꒯2���_|2D�4.��߼3�����.�[�n�7�������s�]��Wb�M=��P�,�S	d�C�)��ι�qcbܿK���C-�l��� Z����2�}m�J��m���05�7�{�Q�s���4�ߡ�V3/0\�����:�֞�9�����l�*��*H���e�O���v�Ye�^� ���IB܁�"�Rr���M-�[Q#��-1\W��^#C�a�_�?����-�[��Y�6���	���%�v�%��rGHv�C𢬶��5�\J��S��U�n O��P�R̾�1���?�P{G�G��>xZNd��0����e��DБ׿@5�	�)5�4���O")o���>�����IŖL����5r��&���Q�	���~���������&���F.)�QX�"����6J2&5�����Xl��,����&6����^�n(�=�7bl��9�n����0��:
��?���e*YxjS��9"]�
{#�rq���	WH�%7;"���lތ��S1�������S�i��e;=xbF�'c,��}�(L��lI���  c�) ��׾,�v]/]��7Gn��P�;�>$0K�"�ܮ%/3�\�=��`�N��*��������J�Ct0��A���U������B�r��y��ֳ\���J�-Sן�~����M?ő��-Yyj1Y��#�c��}��lu<8.b�>k�W�w������C6;~���
�(P7}y9A��r�/����UbvƾKo���}}��������h�xp4���0�+K�ۻ*�L�\σ-���,��p6���}��:�2��&��X�G_4ڲ�33�2���~*��^�Y���Ӹyo�)0c���x �D�ҕw?�sol�W��p�+���1{�P�BSR��h��>�2����_��㐐z��s2�2�����@>��6�b�������mE��-fH��Ο�gU�v�$/����g���͎�zQ��E���)77*�s�*D�`�jyc;X�����NvÅ�]��F��Z��ᧂOE��7I�TO�ό�ﴄ�-Q@�qt�(�]޽H�a�!��AS��%$�J/p��Aׄ��Bt�Б#H�&ԏ܄�J�pͱ4��w(Mg�o?�S��(ƝkzI�ü_��ʝ�𮀻�S�Ö��+�I~<��U�v�����۷ x��Tt`>�U�	���~�����{�r�����h�!lPf��;}��	�^Ma'��� Ԩ���p�|%Ke��u@~�>��<�}4﬚���
0Is�<PDN��7��a��֕�:��x� ���*�o`B`� �Y�)P6(	}3S٘�����&T¤1�G!�s��pG��Ϭ���}�H͚�Nr��݋�~�˥�k[��~��څˮ�%��'��9%�Vq:��T[�#
�x°|r�.tٯa�w��s��<]��۽�Q�����ۛޝ��Ӗ�~�=oy�՝y)Ug�n����R��Ec��h�v^�\Z���n�lJ��H�3[}��x�k]>ʚ�J� u��P�ɟˢ0��������4#kB��FV#fe�ᩫ�j=O����ՅF<\�E��u��yr$�΀�7_2���D�k3��׳W��2�Z�e�-o�(�n����3�I\�pЈb�����^��q.$W��<�}j�һ~���0�κ���D�W�!�@��4�+�P$+��t�ȼ}Rp)�_�}��{�5��L0�i��r��!���Jb�t�gwfLYT�n>��2�R3�������=	�qh�2?�ua��
94)��OZ��V�	G~��G3�-7�Z}3t=��vN����z3��Ń�t�g�>v#z%^\iu������O-*_��t��;�/�����=�'
`tm�]t�cy6$5�5ѝ�JaIa��@u^��W�Kp�D�R���<RA���=�㸅�ry��4��Q\��=�_�,�g%�]ǆ��)-�3H����[/��¬��)ꛫ��<5���\�_��.Z�T�5���!�vP������b�������ø�/"��A=��ڶSaP��)F|���m���|R�b2���������
�k�k���9AR1&wu���5
��ޖ1LY�/��3�ʦ��!����g�a�N�C�^�D �P���
%>ƍ�xe k�!� �q��z9},����K�R��b!V�� @~"'d$��JL{yIW���D��P{��ӣf	NO��6��Ds5Fr�l�E �q�Js�:#�7�����uF�D��WWu����n�<��E��ؔ7���t�
Z!�xA�,�S�~��֌�_�0����M��3���r�	]$�Y?���`�=��X��ˆ
�	k�Lq�TQ���y���+�,�4/4B�����CZ2s��H����f5Y��|z=�����րSL{!�Z'�����a��� /T$�8F��¯���,��4�
�=*ͬ��iJ:�V���O�	�'N~/�����S��GzN��"%�fo����s�g��4a:�0L�lL�w1h����w�{%q�����u����sՒ��nUH�p�"����*�ё��0\��wv�M�8��/���P�{E�uՕ�A|�Bf��O�P`���E)����9�ý�9�`�zk�t#�Š�o9+�9�ҝ���o��G����l�G��k���F<�Y�)a���#B��ȥO��Z��O�R�9$�rW���dj����z�����&Q���$��vټ������_����Fۦ.�l���l�]
C�Wboe�ޙ�]�tLY���\���v1ڬZ�@��a���Ji�2�NJ��Z|`*G� V��H��)6w_n��	��[|���_u�68^�>�3�N���G��/N��U��'�1�҄������!�������ķ��߭>=_���\Ë⍧j�Tt �0���AB���	d��8��q�4��H�����#5x
�:�����t6ؘ1S���f���9t�l�Ԝ���7S(���4��wV�ڂ�G��Э�c�����s=)�W����z��CiLԄ�D��OMAN�!P_o����̪�$M�!�Z���gVE׮D=��Go�Fʼ��Ɵ4I���1�-`�G�@$��le�D��^��]��_�;ʳU�HPAMC*���x���S��[��A!��ۗ�>O%Bjs���Q�PP4a����E�X�n$�p� ��`4��Yf�)�c2cN,93A�+wpյ�wΙ�U�'������zc�f\����i�����YA!(! dIqՎ$����$e���E�˴�	Qq�y��3`�� ��&/b#���}�ͅT���Pl���5V�2$J�(CXZP��z��|)�?���6Ϛ�Yv��[��v5O�l�¥�ͬv��#*��G�ma��ϊ���ׅ
�vH�B`�+b������AF�C*}��
giH�%6��o�'��ӄv�r�G�� �F����#W�|"�����!�U��������rkh�֪�4v����rw����!TDCp����n3�,�cc_i޺i/�*P�V"7��\Kgd-�m
���F�J`�.!��0���QC\%�볈�%_� �T5�f�+�{ot
cF���]��Iz2ڈ4����u��~.�}�&�t�e|aO�Z��[	�����{�P��7)ѱ��j/��V���5�I��ʬT���K�	.�߱e7z��~yVF	��Ҥ%�:�n��X╦g8$:���yG=�	��7�{a�ԃ��9��gw�z4n��2�"]zq���)%���4Ն�*bƦ�g��-��B�.Y���XI�>�"�r� @F���Ȓ?(ˡn#�͠3���3�D�+�]�M�E *���:�]ڠ�c�:9a�@шIW�ON߉?q�&ne��?�{��$���������Xu�a�p�>���Y�an�M�(��1;(lo6i�yL���w<�/��勒]熎 ���<�^���ܸ;�(����8��BɈ�WD3*��m���F�ffp`�!1w��?��#�f�}S�5����G=-%�cɤ~o 
~Y���g�گ��;�ܥ[@-�ۋ>�z�ف W����q���A�
ܛ%��I��;�ұ�O^����#��UՐcyk�2p��>�997�^츿�%��T
�Yͬ����g}���Uv\�gq|�\R��Qdy%U��"�5�+x��<qAǏ�e�#֗�|�E��=y<�䑫t�+�y�J��g�/�ˏ*$:Y���kY�� 5���6LyE$�	=�2�̖\��6z����U*�8��Ml3������Y�J�#\�)�d�?l+ӣ���k���{���9��Q�B�~�W�c;�\/(69�g���� ��D�A�;:Izȍ��E�Y��%��܂G	�_z*a��ʧ��A�<z��骲�m�

1�����#�W��	���$�eJy�LTQ/�os��wd=�OJ��}���k��uA�h a9�訠3��!w#���ߑ.�[��ŚMp������$a�JӸD�NX3Cб6HW�E��jӾ~���jl(�E& �8\=j�mN��@y40���q