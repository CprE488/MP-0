XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%�M��P�$L'%�1ju�\d4d��JO��V�Ybu9�<:���^@:0���Țg�=ȧ�A�p��:�݊�2œ�|mw�ePy��������4���Mxn4�m�K��~a/�X�}��!a@�qdz�!�
[���L�ia�84C��?L��,�,�m6sU5�SC1�#,L�g�M���/������?�Ӹ���^y:G�uX���<��%���,cy~����JV��;9����=��	����P��x:&}��=B����m_�,��M�j,Zi8M�x#�|�^] g�A�����K�o,jm���6ɺ�7���*���)�Vկ5CW��d�csV��v/�Va�cK[�����kgh�6���������%�w�wm=k'+�+�Vs64?oL�f[Dц9�f�j���r�2+�ʑӤ^7���{e���y�]���b�����hHƩ�cw�F�M3�Q!%��J��l��&�e�Me���� (�S�ؕ��G&_���T~�����f����4r��)w�Z2�Z��8�Y���Dݶ�3���^z	�:L�Mܝi���|��2�xp7J�X����%s� ߦ��]0Ղ��⧖X���7�nq1u$�[r4�Q�$g �B'�l�/I�o2+ř�uoL��~}���1��Gt�b?m,����M��j<�����S�\z����ȓ��ٺ3�ƌ� <0������аD����J6��y�.��8"EUd�Ţct����&��޼$XlxVHYEB    3fdc    1160d]ј����[�vj&_в�CxI�叅�ŉ�̯8B�\��_�X��e3KuS�m��.ޡ�Ā!X�m%�[v��C�^T6�#&E�ۦ�o�\%2�q����p|Mas��q辨v2��L1���
�44ΔpE�g�||�B5	0�DB0�D��g/����yd8T9-�������r1�=��D��|7�C�P�� �[$�F9s�����i��|���P�� o#U� �\E��*j��N?W�J�
�w��ږ0�Z��/�g�S��xV5�/�g-lD��g���Т$���A�햎v�׹}5���ǝ%[�đ��خU=awW�)syݲ��9��40a�٨��3�f��e���������p5<�D���4'�-�^He1��裉P,#�����Vh&�N���hd�{�>z�\(��w.��a�*�L���H���vq�b'�#|�D&����<�&�*��0~��ke�ʿ�3@��؍!'�'̈�QIp�-��*�{��8CA94Uv�YP�ܺ��%ѡ 7ܽ�58DC��H����c���8�壇_�D�����:[�쌓�n�MIq�����ߤ�_�O�n��5XN�uH�&��O�#�z��n�Kb��'[�������:�
�<��=��=�!m�_@����⺝��	��7�RV���/C��[
ۥ�
!_�н >~��Ջ)M�"�;�ĸ7�Ȍӡ�^7��W�c,��O��t[$ߠ���rd��8��/��,��s*���y>������đ�����笧��� S^�\����|X�У��c��\�|j��W�%��t�@��U���L�2'�(��Q�������`�O�z�5NtvyD!2���6�W����������#�9c.��m� ��Mw��T�+ê�Pߎ���1A
���*�d��{��a�z�?��˔�����}�rQ4��vC�e�z��2*	n�\�摚3�����t�f\)��גw�{4;��~��
�����L��"���6 ��Î�SI��3Xbȥ(1������vޛOO����%���m$ ��/r����*��3&By$/����%���xB%��|F��O��Z�z`�N�;^J�<ǥf4��ٲ�K�fO|�7��Kًۏ��=�B�h��W��]�(퐣����N�]h��_
��;OyaY��c)`��2��ŭ~�"�oɇ���tt
�G)��z3�J1���N�WA^�LP&+��W�2<�����PW����62�5&�8�fi^jǡ���2)O�˄zc�$��]��=^�(����ƿ2(ad��Dɠv#a�|<;�Y��86��{r��������8��}xd����S|?N�횯�%Ep���A
�%�|�ͬ���	�Ý-��F{� �7X���{i ��Pr�ݍG�TL���-E#���ԎL|��F^��� c���.��?��  K��8S[�����;�gױ�:�U)a8�M�����ֶ-I�ph(b�ZZ��$��Q�{c�},�����ó��Sf7��qR�&-���C'*��Q/�bZ��M �+�K:. I�jP<��e���1l��:x�aKp���֭�P�pB�?����4���^
	(�&�����!`�B�'ų�VK�1��D��=�TdcX�3���C�����|�l��t߿���IT�q�jͺ�ܫW\�|�� ;�*I"M�c��=@������kd��$}�2���K�OVW�p�����ĊlesS��;�'����{/i>���6�lHŴ9Al���?�a�8��)倵w�����U�\�l�1�G�.�G�u0*h��f`�NCξ�:*��J�	��V՝���	�1���+5��76��K������|Z�=��"b�����.J�-�#�u� ���ޱS�%W�hZ%Lor��L*���f��<��
O���9�ġ,�#fQFz(�*-��d�2:�1�Y��A��.��=�Z-�\x���Ҋ�k9n��*\J��_�}�9�P�k�
4���T�IQоa�B;AvIb�4�C�ryW�2T���ߌ����4�M+�f���0r^�'�Ϯ��[�>�ۯD����F�'�8� #���ք��P�g�g3��V���m,��d�qCx���s��>d�-aً[�a~�￟�6����~|�v4'�裴#�}��U$�Q�`���W��7��]<�|������ �����%��(A��{��ڒ�\�^������7��b��+!��r�W��$�o��\˿:��P���^̦o������IX2�5�eY�v��Y��OU��7$�I[�S�@�9��U����rw�=m�.���]\@Juፗ�I;�N&&�.
W|dV��8�e�VUU�؅�!������yǦ�
�g�C!}E�[����K+�y�?�-�t�x���ɢ�g���:�SVx��
�Ԗ�]0d;L{��۰Z��>m1K���+�5��3��Ŷ�5^���`ߪ�,���O���1c1&[}G�f��F2Uu�)C�{�Q��d>���|����9A��ZP���i�Bz&i���\.6���?��.)�l��y���g�'Wc5� �D=�s�m���$��DjDo�)������S�#��S��^S��l��Ĵ�չ�"������,W^�����*~�V�.���5>��ĂÕń@��ʛ�$y�'����?䕳��5JL��(g��mg�Z4���B�/�tq��7�Ud�gȁ��r%�S�SyѤ�=���ژM�
�Jݞ�ټ��|e�pA��	������S�E*Ul?
 IM�c�x)<E�����ɕ�L��������]���!S���W�Dr�Ƨ�ꊏ���-&�/
E�#ZK7m<���oɦ�)�Q(�k�mPN�����W �r��T��Ld���{���^U�'��</yr]7V������,5�L6yǚ�/�1o$b6Q�;mǺ�X>�ɨ��}]3�p��8�5Z$��� �����XNx�qv���N���a"K9�O����U[g"�-��`���Y;C���ν�h L���l�9�m��f*��dlfg�����_�s��B!\�u���{�$��]��QM��Q̐#�R+س��;�����YĹ3EM)OLEŻ�x�Hy��P�h8Z��uv��q��>�?��,��[蠗����z(笈4#�p�Ћ�3�G����3�P������+Nb�(�(x����M����c���4� �ƏdDz"�&���$��AK=��w}Q.>B�M��8���
��a��F_G�:��@�r�GrA����l��p���\�%/(/Ü&��R_�Ѐ�Z�>��bC
ݣ��D���g7��f��qCwa8�l�䄣R�r�X��;�4���ɣ�b�5�b���B.�h��w3�9�/l)���z�򢻸o�7ĉ�'��J'��	���/������߻^T]�u�}��[�*
I�6܋���2�Ʉ޲B����D��Y�LPؔ�Ή�.;f?�J���ͥ�I���>����XBA���6��ˎW��f�cUL��D���]=����H�_��N����d��=r�N�j`���Ƽ��\}pbѾ�����'�Q\��h�䞛��,u�8#�c98`���y������6��<�k�7B���<��&i8����I��ǐ��.w��ĈGUD\{\~&i��p|��`�8NB4P����R�.x�Ռ�{|~�d� _-����`<I^��3Xڗ/�����;9�����d��4����t#ZG0��۲��fm�Hѫ�z�@�/���:N�s��E����I�3O/4�#��5ܮ5�.8�2�_/�:��J�0䲺���ˍ�3���_U���7cT��o}�4�U�t�<����W�y½�щ������Ճp�����T�r�1e��9�M�R�f=ߜ�g�H�ڤh�p�""���e��)Tr��9�
�/υ�ƣl��IC�|��9=4H}�g�պdT��0g�]/�h�s������c�����O{#����kD�M��xe������C�3����s,?�=��?� �\%�I�$fy��s^n�,ϏQG�,���
ܒ���Jl������z��B����r}��q�HSW��}Q�gy����3t��"e�_��2Q!��Eʉ�F��w�v�1��P8(�˥!n�����	=|n�[/�O�I�o"2�`eVP� Zza �ٯ��J�ǣV� �����s 4/���}�]֡�w'�K���d�����������v�=�Q��L�@5`�4Cc�Sh�3�z�m���ns]G�ɢ���#�������Q ��D�
Bk�j.!m}�ɠ�