XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���S��F���6���%x�Q�gOHxXv=���C�%`}���/Em�;�H1�q��U�Oh<eU��n�c'�9w=h{�+�4.���#CTϛ%͓������8mf)�1��C��~R������Jyѹ(�O$0�3��Q������/+6�s�M�;������"�����;���Dj8&W�Z]浠ILb6(.�ѻ�b��A�zu	ƒH�w:��\���� �=_����Ahc�t�1'~s$���D�ܖd陣|8��u�(��2�9ݰ?)�X�8%w��n���I�^�+ԫ7?�6��M�f���W�Iqcl͐���Pc�r0�!8*�2a�>��>�g��bW`�
A�����*�ݖQ�����?�³��"��L�q��3�Ƀ)P3)阆=[&@��c�.�,��f|�;�
0g{y�Y4jց�C�M���������Ǔl�j�y���vv�M8j���0��K7p���R�yowWA7��䷚��ٞ�=�Rkρ��ua�T0H�9LL�}���{�Y�y\�{)��'+���s��P�iEqwu��u����J�0(24h|1�r����Ps�ϤI�6�Au��W	���ԔS�#�j��1�1����7`�e���kY��/�_�ⷷ2��.�?O�{0��4����R���ې	n2�+������oX����H�N�žj��X�����j)׾n2�>�$� ����1^|�q��Q[3��$	0��G��r~c?.��q'�#��I�{�G|u��XlxVHYEB     f6d     6f0�䗏oX4Ÿm���#8a�MZ���5D�!�+�F��� :
�Ԓ�O��8^��Heƌ�����Œ=c��m+K�V�-7�&��Dy��asu4&��3	�=(-��7��fe��R�b��+�d
��k�+OJU.DGX�������K�W�qO?o��LN�O_�?�/-Q�(@�_��7�d$Hk!{u�)Q��a�Pr�y_���Pp|+�9�uu�F<R����χ�����g�.t~޻�A��n�Bn�6�4 WWDf������aR�;$��w������o�'�foK��]|wp���l�f�V��%2%���Z_v�����w��-<��r���J>شB�mN���ΰ�\��Lo��<̧�xc��6+ߣX���ڞ��q�{x<�E�� 4��K�p��Vaf�	$ɠ���m��m�+X/|OQ8�g|d�oN�8���2���?}[��Gm���}7p�JK��"��A���GOR�7����H�L�yZ&ܜ�8�E�"3U����x[{X��%ټ;��/k��xF���n4�έFvĬl���$w���k�ZA0#�|3���a+ې$��{qu�������BPe5O�\�݆���t��D2��ɟ���.v�.F���5����(��-� O�s_��X�"��n/�gՊ�����"I%Nm���I�,��=�|�	l��5� �>ŵ@_Y�b=p�uи������ULC�y}���U�HyX}�_��|C��1;E�|��]��^���I�eا��>���W�#��kJŦ�!I�n�����%��&y�NT%�''bܛ�<N����gs��!�pl��rs�u� dڿ��-�sZ��:m�&�i$$�kp�(Q6�-w+�ekG/m��|����+�coqG��V|��i{�;��Ͻ	���sl�qR�1�T��Q��f#�'^׃�~],M-3�;Q!]v�� ���gKXp��c1ו����W����,9s�����X�N�E7`}[&p��M¸q���x
eu��wK�{�J����N��̊���rS��NC]��+^D�0@m���丏�]��Z�jD�0��{Iy<Cr����Ov�r'�K�� �ۉ�c�ߔ?�X�go�0�m4jONU�`��ց27`����~��kW֦֗��۳0wg��v�Z�����$���6ݭ���5n�̙��(g����_�O���Dj#��v��3e������z32p�Pl"�j��U��1���Ц~�LK��2��Z��CH{� ;חL�C�̭[��k���ʣz����J&���Ř�d0G�\{�q��3�&L@F�Q�]� H�S�@�� d�>ddw����ܟl�˳r�;δ��A��W���q�`e�kY�5���U�ķ*TgײN�-�����@H#[���g���K>��;W�4������c������3���sb�1�CCYR��W�p�m�b
��B(Zt*8����Q�ͯx�U-j�-PH�i^����X��8�:�ۏƎBZ'g����i謊�Ӹ�߶��X��1��Ց�~h�%�����L�z{�h�򀥓m���*��&��ɯ��W��5��
�u�"1L�%iS�2<���e���]��\�If�):�SPyˬ�_A�Ř==����B��&%���2Ѭ�~}5�f�>�W�rm����|U��6^���U�#g�Ab�j���f����(L��*7a7nK5���V�(�^{�l���a�Y}�v�0p6x/Zs���e搆f���TEb�]��@