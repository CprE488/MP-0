XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����`x,ўkS����I��4~�	�;6��'�zq7��?����4�*��<y��akzy�`�1�r��'Ib�B�@�	,6\���*��Ӳ�,G#|�mU�%� ĂmE��
���形��Crt��͇
���kn���TPT��y���^L4l��屡���W6�QK��So�'�UJ3x	��@�}:5�Z����dN�,М���f�@g7�P�kQĭO Q�a,b��+~NU���0��V��9����&?ueBo�����
GYF�8R}mv��)�u��e���Bx`+�g[甴��O��<���>�q@6K�����z,��#@��W� ��+�"��:���Ҡr'=kp�Պ�N�N�?�����Yc,_Э�D�M\o��zB ��%)&.�Kt���o�=k��L�ײ	��c=�~΃��%#��N����I8���/����
sc_*��	Vγ��׉V#i�N��u|�W'EpA9|��@�vGk�.O�̰��)\	C��-n���%�9� �t�
��Yd�_zԛ�L	3
q�PV5vf�????�qt���.�����F=Kz������6��V���R�tk����P�D6j�g�+�Y��"y��7yi����N��aڋ^�,4],��Qwϲ��y�W9H���R��ܨ��fA�Yg�p=!)ɫnna�Yi+�
�q���.N5n�w�O;|{X��@~�|�z;��u;�C�q��3
��(��n����&vd
�Du��"�<�%B"v��0�%pT�T$�!�XlxVHYEB    6014    1840^@��wx�*z�ɍ w�^��L�=��q�'��2*���N�����/PB�=�fm4�]G���Ib'( ച>t����~u?�y�~��M�M֬?�L��M�i��Q�:���PQ�-��1�	Л"��nE���GzL]D
eڂ���8�>/�n@��_�n�/\��,��e�:�B��S�lK~<�D�J7�X'���+��~c�Q,GF7���AY�[�rA�ְ��>
�ߞ����a�°F��zB6������M���x��{�aq���$ ��}!���C���ɭ�S��N����I�)����<�!Y�s��I� L�F�>�>�'-9���Z_���K��*��yl�0�Ek��T$�v5A��S=��r������~q��HW�(\ y�N���G!�L+�!�a�׉�S<}W���=$v"�-��y�X�G]��Ѳ�]�|��������ۈ���/Ǿ�y�o�`��`���K穁
�r��vSC����H��g�]�fe�;c(����Hg1+6�p�����g����y0)*ؓW_%_���&i�U��ю5�[���#�kD�!�Q�k��,�#}V�\$ڲ��O���bM����&����V��T)D %	,��K����'���ˎ�u^5+٪K����z��`LZ��E�9�P���fEP�XE�� �CN�l��s�p�LC&4�B���FֶM:$t}n��1i[�\J8-ϹPoIa��-t��@�Q��yឍu�}ő2���v5L�_Έ灐D�~0^����e/�%e�B�k���!��;�Qo��s��Y��O��뜆�,��e�������j�G,G�{�G�Cw_�v�?��%x":$%� �v�޲��)����ePdj� }��8���q��Y�)�w��\���}-n8!OB��!�-獓���TBC���h@b��+^����"���w� l�"D��/F#���پd:/G9疂{��3�%l�;)N94����K��v)��W�58;%O]�Z	��%�D*���P����dT��{3ەG�Z��lL)H7զHa$��|X� ����ҨI��^#\;KQ�B;��h�tȳ�5�-϶w2M��Z/���]j�C�Ct'�{����{ϫ0���Hb�mV��6����i�n+ur���[�?���D�ۂx�(É�21Fj�� ڂ�G*5�k�7��V_�lw(��W@v��d@�{�<�*� <����B�`��$'l��A�u�@�7W�x�:m�����Q)S�ʁ<cW��N��vML^�/��_N��N!�3Gq&y�W�4��~ԕ�n��L#�CY�o'$ԭK�w�W`HJ���G_��}��<�W��q��I~��c<��X#�)�@%P+�ҡsɃJF��mA��KA��e�O�=`�R$'lOϭ6]/�0��@��.N��*4�����<3J�jg+��1!)䣄c�ѫ�Vx�.�ߩf�C�4���"l� M��>#Z�.~*�,��*�f<���
;�$��n�9������S8u��"<f�=��-IJ�T�2.�dņ�6G��|j�-�!�*v=�i�G��}����gq}l\���	N�,7�1-=�vs;���G@u+"�"��J�Z�Nk��edM��,m_rR�t���0f�'*m`���o�(C�"��A#���p�v���Y���p<}q&*�'�9��3OY.�ڲ`|����o�>��(�������+&���=`�U8��#�j�]5s��;]$¤urտ2Rc���GՆ� ��_o�Ʈ#�V���#��E2���_ad�a���t?�sb�Mvb�Ǝ�9M�X�u����g:��9���@��X �:�a�I�����9��� v��T`v�]��uD���bJF�xe؈#���@��$�WV5��Q�g`�Y|'K��LY} �	��9��s�Y?�Z��S�F�L�X�D'�n[ f���^.��2�[<W\��\7s���8Q��W��7��q�:��p����3H���^�5��S�PF�ڃ�>kԶ��e�za�� ��^d�`'�]�y�	�P��YdѺ������znݸϺ��]��|��=�P1tt�_�C&�8f�*�ٯ�}=_��a&I���,o]���A �7���0ah���lC��r#��*i�3!���[;�o�����{�x����G�� �r�7�Op������L&���J��̍�u~����[j���ћ4^&���CP7S�M�EuN�ԋ��Q�r{����S�%�j��}��_�␞���j���Yi
x����Rz�φ�438���jz\g�F`��rJ�Y�߇V]��c��g�|tM|�� >/�6�5�e��Qص9Ca�0f4O�j�W�� ��f�=dV�΂;����|A�bl/���"p0�E�z�}�<V¾��1��v�%�nH� g���P��A�8,�3�&'�!�M2A~B���Oh�2c��r����`Y�xL�Α����sܧ��Y5����n�
�����I�x�H�,��D�HB���؎�]�y�4��� ����E�|�n�U�
�?e
┿w��:�G��e�f/�M�=��+���j,���fې	R����BNi�4��Ӏ���Zl|��n�|�Ϸ��~�������)�L��i�8EB�u�XL%�}������nQ٢�Ԩ!��0�>�Z+�ߨ{:����6�I+��BmgX���u���4��7Y�+�I�Lz!J{��e�'jcaynd 5�b	�C�W�r���u��r)Ll��%�T�
~��T��m0r3�\����B���$X�qP�\�Ta�<ƩM�zn����ڨyѩ�E��]F��VQ�%�;*[E�!���@�c�J���f���A�մ��Aӕ��k@�L��R�۱�qw'3��e�Y��oaJ�f��'^?%�V)��<��ιs)z�Oi���ml V�
��]�����"��5�_n�NjI��Y�w���T��.�3M�	�e�]^��2�q=�v��%hV�Tʾ�b�Ì_&{C��ϊ�|<O�S�	;������!���ۏ1,7M��H'D�Z|� �"�^����=�T���Jv>5�1�sa�.��S�I�3���F�a��_�2��� !pk�jk�j�R�z0�u!��b���;L?��
%,O�@ɐZ8��p���]��Y�]^Ta�LT��N���?c�ɺ�����_����A�Q51@M���V�����Լ�̓r
-FR7|ܡ���ؕw�Yw�ʬ<`v2���h	pI�ac���+�Q�i�>q��'�:0�v:��V�xS�Yïʮ����O:-��U�,y@��pow{�J����LHy|���Z�H���<�;�i!�@7����Y������Μ͌��1j�){�5�Q�MfL>Q��_T�5�G]�B}KP�U�G��8���jl�tkZ�e���2�|�p�tv���5�E3g�n �����;�Ee�>`����� �1=�d̟#~%�t4#�����;Y���d�:�?3���)y�����8}������'pJT����g���Ѭ<_�ڣX8F3���(y�8c�w��=�xl��D���D�}|�m�����~e�/ȱ)�>mĜ�&���̎��{�,�%�%��Ҋ�Ȃ[�sb�D��ȟʀ[�>�C�&�^!���e������:�QxF�}�ʑ�T4�5��7�#Ϳ�'�L�P��<{/�ު�)�n�G
=��v
��{��/�iIй�y�Ŕ�FUX����=�<�]��t	�w{f��쓼\�,��s����'� :g���E�V&�=��&��;>nKQ���m��UNF	rɶ�X�Y��^]=�|��ٍ ;
y0�xg`�YX\ڲ}U��>=u���!"Ci�g�m.u�[v��}�x���!��f5y�j��.`�`��w����|绸l�Y���b�Dao
8%X��L�&����x�Hw�G��<�&/�$))����qd�s]3�����H��yOeC�9��g���\T �^:�53!+�1��e�
L&K�3O�X5h�\�7�����"�G?��Ȭ��9x�!�\���YJgE�U:��`%�p��u�0쵒�	&%6��ٸ%c�T�S%�ZVo�1?�Sx��S�b-�E��e�Ҧ��65C���t�����y[au�ԗd)]��K��q׋����s�m�l(@�=ę/PÚ~K�MP�����{4��&�}�ӋB�� ���=�#���Z�s]�ygv^kˋ�͒���?nzx�=�ø�dօ��(2QV��@T�F�˂�~x\�o�g=��n-w�>b����aV"��H�5�R���#�����zT�� �J
�(�N�|䭈�R�1�L�x-8����pc��+�X�§������]�6�.�{����v�&g�k5āB����M��¥��oz��â[�N(*�T��<�������#�"��6WS�8u�;��� �����S���T��>��?~)7Ԁ���&u$=��L_��R���Q�a{8;x���K��k�,����l��D�7����a�A��#GE�鱎�)��Q�9,r�8��K7��a���p�ĻB����6љ��#V�L��_��>�gg-�k�"�7�yv2���`�~ZA&E�c�:��sy�j_*�wYT�a��A(Y�p��-E��7�w;*�(bw�lS��o+��a��99���҄�}��IG��6| �OF���t�l���e'�Iշ�@�Ŷ꠪�P٠�e��a<�TK�Aײ����=�!��,�n�w���$M��a*^+������kv���?��$�0x8,�WTN��>��VXJ�d4�0�&�����}։N���K�?��H��_��u:ԑV�	_�.9�^_�V��o��a{�|��i{����9�ك��*7liz+j� d&��;we��Sn,�b\=ڧ��P�]*�C3�ￗ�Q�`�H�~���I����´����)&�.����Q�=�ï�h�96��Q��1�&9�H�s�xPDڷ� ���Q�	8z���9a{-<�U>v��us��pl��������
\�u��+����L!�rfZ}�]�p�����q׶�pL!A��L���R�9�$�Y������z�&�Z�������/�>�`c�L5#m��~,V�g��8����q��*[�6�����
9+w��n��JZ,`g�r����૚-�E�E�$�!����D���Ex�{#����缝=������kȖ�-�Rǲծ/���GO�1�L��7,�sb�L"
�����|��ge���j��U�"[���N��⍣��ڰ���«s����n��F-�Aؤ70��p3y8P[�%Fv6��}p�>|�Q��D�Б�H�]>���씕ɩ 8� �"@������G�\�<G⑭��m�a���G|7"�w���|���-ԯ�a�2��B>�+�|�m1=7�ˌl�2�P
�__t�ن��B�N-�?:��O��4�.����Rq��>-�����Z���LW�8�dWf{ڵ�@�R��X�2�Kʜ���{no���`7VF���b��&LϾ �k<�����e�
�*NV �BNG9<����εF������S���f��3�D͓fq��Z���#��;�Q!i���{հ~�)�bq����c���ap'2��Mh$�����@��:	�b@ۭB�4�#����x���;���P�"���-b����c����R����JO*��cDPL��_��	1*�� /	 ��|�D��I/{�� ���0��,�w�Y�AK��(0l�G	[���������
D:��� c��!��E���c�?�p�p������ޓ6�[ئ�t��qFjW�6l~�|�\B�11�)U��'�����F[Y�����y/���!��;��C�"��Y�ab��y�E�f,(�:4x]!��U6s9׋q�!��(K<�C/�Y��mf�n�,�c%&�P��:�����MowN��o�����>�a�0삵�+�F%׾x�V�<=�R��P�y�r
uKxA�82����BB��2�