XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&a9D�D%�����~�E��~z�Z�ڋ2�%a�8�g,��c�zc��-�����y�3
o����^�ְ�Z�u�P�!��b���;as��݊�;��-�[��̟T2���!9��T��?u����+jl�׵�rc�׃�e��>MY1\��I
Xi�ō;	}���g5�;�>}[�m��+�ݛ@�H����9���6��A��1�x(OBpK��s�c� I��sh�V�/X���:RD�ʨ��d�w}g����*����x���K-f������>t� ���1�_
�
{G�em�j��"�+8�$�W(f��T��)���D��?'������zdb�)v�7�{,,��T>�x �E}t>?��X���<!��@ڂ2t-.���IH�>=256Ӥ�9i�L���8G
�(?j<a�$�Ȼe�"����h��qDl�:W�s�{w�z��93b�v�y�e���B=� y��W"��,h�(G-~%X�Ay=�����w�;�UP�?�hMᘕ����)/Z�:�[3M��C}X��P��Q���/Cc�A_�|Ȱ�D���ЀO,ݶ-��ކ��i�z�c0�$�[J>;�by�)N�+��p�]QP� ��v^�(w��ꢧ����^�_� ��N-	c,��B�&PF�uP�W�4�C��D����8�\��J炪��Nq}���)����N���%^��d�>/U`�ц�9+8g�n�+K�)>���ޢXlxVHYEB    95d3    18d0�=�GU���߄���O�Ƙ�V"_��%<�	ŀ�
��!0R�[�D� 
"�p�,Ϳ��\�$�l�M������.m)�=_1*gs ?�S������c�b�)"�R�K� �ֺ��l!����F)��h��@0�������bQ�g�����sЊ+�IZO��ݕ�Iha�@48�Gim���HZN�>]�������� 5�����8�ro��82�9�M?�|�����~(�^�Ӊ�5���F�%<�-N���U@24��aI�o��I�rܫbc�YͲV���o5u�m��c�:F�����%9f��ݠ��3�6H�و��������_iJ�ͫ��j��nS����c}�!|ucT?2��5\!͡�����t8��܊`!�h�#�I�G��j�/�!''h#f`�X�#����ɂd�W���5�٢�q�h�(��`�.�ho��ٷ�]80Hw3�� (oa����~y�fY<Q;��ݎ��,�%M|�qM5���k���L�L1�+�`2�2��d��._ة_lL��p.��1��#Ź�_����U�w��6c�G}��M�Ga��W� +�j����-8�\D�aG;&��,W�THq����~z��v69coW�����;5�vDᵞ�9����-ޘ�Hg�/�i���������>KdΧa;$��:��T(�dF�d ;gi�Ěp+�!N:#D�O�f`��h�L���}c�� ��c�]�Ƅޗj�e�I#5�l���_���M�N��er�&�v��VW���3��V�^�OO�/�3�v�+��Z�	��ߓ:�`�����r�?V̄���Me4a�4i��0�&���t�U$��>1�>P��?>�J�C��Y�f�}zYa�x'�5*��!R��RY���n~�ɍI91|��\��d�5,<y}�,v� &�^�lgm��7?3B<��'e�	�rܠ�K��?���7�����9�QQ3Ų%%ˢ�"?O�������j)$��l�!*����8ԕ��t=(�	��סq���o�N�;�Y!���B<���m��R��Ҍ�t��1�O�$�ǻ�>�h�;��^��w2��,\E�%�w���>3���s����(�Ve�_� �4W>���'o����D��75���V��WF� ��	X�9K"���A�mWE�gXc	�V���Ģ���L����S�x}0d1���Tiu�O�E9�� ���F�[����/I>��n!�1lsQk{�zO��)��a ��S�I�?�x .�u1�ӂM�E�Q>ԑ*�zv�o���R�����У)��s:htȥ4u�P]�M^�&�p�<�Z��orSJG��fpKo�����.?<��������c�@<�Ψ����I`K��a"�P�)��;U���i�ښG�N�2C<��.�ڹˠ�^��vhE���g2���HS`B��_�7�¼�jij��E`�@�vK�15���e��lꤑ��̟���h;KF��U��v�cͽii|3j��'�l��@7�'S96}�݀����O_�H�l�&�V�8�~זu���ϵ��s
)�c�+T�Mcp��&D8{�C�J<Ktm(�e<�+ΓD��M?�_	��$��IG�������,���WK�MhؑU�b����l�L��*f�tA^���Z
�<X��t#�JQ�zc���^�$k�:�;:,d�"'�����~�$�T�vDf�RE1f�9/y�]`oޓ��c�x`����MDnհ���{��X�{��š8�Kj>�T�Weyg"�AL��JY��c&��z�fn�[���s�А����`9�'�-���4���#���V���<u��������m��6)Y2I������ߜ_�d�m'f3X�;�Z�Y��y������#��h�}0A-�]��J�|�����s<a���,V�N���!�����f�9�ntŁ��O�"�'�[��XA�%�*�t�y�v��@�*Aԕ4sb��Ek!)��<l��λ��H;c8bx�/e+�1TL��O��L�P��.��<^<��3Z��v,�����7����ީ�6C�(L�u���%{/�n�٣���*���W�ӻ<�x�������)H��M;z�A����h1X�_��e1|�;��'��tV�AG|�0�N����p3;����1�^g�Pl7�eX �!9�y���k�]��e\+<�S� ,XKo�Ṽ3���n`��=�og/���A�����\����E�k]DK�ǂ�rb�n��2���M�|�6�A����ZO�>����-���A]ZR0����w7�A��%J��c~dJ����pz�2�9�{qZ������A2P��_H[�a��z��1�Kj.ʇ*�z�^� @���WX��.��&�T�)�$-M2�v�b���w]����a��ΝN���v�.����Ͼ$,�n�a<M�M�:�"|�D �*ΧR%�+�I����ɭۉ��%nI>x�Ș�rk�mb�
�=�ULh'� ��j-�$��;(
��	� �ze;����P�x%��ִP�;O�|~6�j��m������Qe�Xn���0l��j0㐾�����Oj����@YQdF"��E���+���Bh����4�V�e�"��.����P��7��[[ïN�:=�L)�ě-Z�f%����'�w���KR�E(�}��kA�dr�ƙ#�׃�t�z1��~���0r�p���۲��nP&���[�tGi�\Ƣ��۽�r79�4�t:RƗ._XDe�s��xޱ�_�ɀW�̅�lC������{��<ϴ��P���+"( ��X&6�>�;�xdͩE��5\��S׻�����l�|�3��=A��8W���C���^ A��W4�I�ŖV��v�ߥ羂�z�4?A�H�k�k*ۻ�Rf�C���,Ɣ6|��p���R�z��A�S�6Wm���a���A�bObUͅf+��8��`�� l­�&,��!��6��o��'�m�����(�'��@�8��{ؠ����]�Ј���=s����@�,�5���#�[�&�b��޳�zI����Dɱj��e��RM��g�|U!(�'�RK��f��N;�D��S�$8v�?Md/T*� �yגk�hƽ��ǆ��a�oJG�K8q�fO¶0C#���4EѪ�Й0�r>R�2��T<�ws�Pi�����s(�@�y]Z0�;�T���ߕ�9lV��D��=ӵ{()�dp��A@'�9�S�Z �i�̢oN����L;":@���Í�M7WyS8N:�Rj�0������☠�&���W���0�P��y����Ao��>����,uk���9�
EG̤\�#������]�:�8tE���2O��}ݣs|��4��/��{�C�[E���B�H_③V�h���rSvtQ�]�F�~b9�5�Z�v;��c�?�>I�{H	����6��-�u��>P�`�^�4�w���N9�ƞ�]�r��6�NIی2��8�z�)���KƏX��)v)-2�����%K8���8ńq�� �So�,=�Q�|\�}F���Kc�w���c��59o�F�'��5�qm��3K	c��ۻ��]���2�7�h�t&_?�bL�N�7>G�7W�Uu_��a�V����)��a���_�8Զ�_'j�b�
��e��0Wjj1������mM��;��A|�����|�(�)Z����-�9
J����S|�(���2
��|aY;�'1s�O�	�����;i�'u��/p���?-��oGO8E�B�zKf��h�-y9[4���m[���
äe�4� �g-�#h�@��bq41 �N�*D�G��$�TӴ���D
��jL^9u_�ϫ�|c�Ԧҥ�1 ��U
�fkS'���n�W1�n(�u�×ΡoI+Iz:�
�D�CF����{��Ƀ7��w�m�" �0�B�L����=�.�(v��d4�y���X%�{�w�i9O�ʭ�er��n�V����;R�����/Y`��`XJ�P%۫�)&����~Ś㘒��R�r����@\��x���`i��<��R���R�2&�,~��ml�uK h�����Hj��G` �\0a��C;��#�MH��fL:��+�z-�3=gX$��~�L�#J�8(������������C����f$Q��0qǹ�Nᩈ_���+h0�5Y3�v�!ėr���C��:��`>�=��R�~���>�F��ɸu�����\����ps�]ȞY]��Ǎw#�*'"�^���|U0� #�p����uI\7����霸{H��g�5��wh&�����z�%�|�0���,B��<OT�D	�S��_%�[>�o5D����Mi*9�t��a�p�ƺU��� ���5^�7̣J�)q{�H01a�@B+D���Ai�B�8P���\�I	�>,1u�l�R�`=�,����f�D�{]p��/�F�[2}	������`��&�({��Q��O��$���h�&���bs@�T�G���ʉ�Y�lP������)��b^�p�D�uT��8����4����׆O5[;�:� `�4���}Q&-QqE���3򴃅�^N{�8>��S�,%�KSR���Ӊ/�^��s�S�=ѳ��	�!����H���G%�HhЯ2�ܪ�<:���Bd��c=��:��F^f̧��`n�� nT�x���Ƴ�������=��j������1���kc&ex������{C0ݮ6V�T��f0�ܤ��d�(>\�=�U�S�gv/��g(w�A\�J)�o�L��:�mT�#��zN\�iX6��2�69���G�X�;w��;d�'4o}���as� �8Q�{�@�9@Ad*���O��+N�n���0�Xڻ=�\�8����(�D|�S�c5.��3��&�����|BN�wG�H��v�MW)���܋b*�^�E�)w^	�<B�s=�2��-q#���P�g;�pUÈ�`u��ʣE׎6�HAu�âS[c�)���l�b����n$�5���砤6^�o��t!�ۂ�Ӟ���/�R9`_��P`+�M�Qd�z�b/�_�v/��,�6�����蹼q��}��7�k6P�\�e�J���x��RУq�����/�y@��7�%]h@��!�sţt<q��Є�}��'0�![�*�{j��U��M�V�#d�F9���}�_d����i:�S��W.��G��#���;�GE����+�&L}@�����v3��hz��g��G3ܛ�Ȣ?��_C#=?�Um	0��hLA���ŀ�4:���tV���F���H&��$�b�RMF�Y ��SL��6�CNEB'g�ro�o����I3ݵ/��Օ�®�;X]{����� 0��M�>���.���]я��8�c��O"@��?�=2���r#�2�O<���x��(`S�U峿D=�&dH�	r�c��2���E�"K�D��š�,-B?��p{#�%6��`$�e ۨȖ�Þ���E9u	�@�h��3��-O�mDiSN�N����:�\��孕^��-�7�J��'v�1Aq�OK�Q�@ˡ8,���A�F��;���p��Ɇ&�o]�PN�6�����%Y�p�El�IB��0Q*A$rE�(*
b3U�T���j�w��������S�хD�E:S�@;�(��T�o��RB!�O(�S��^�����������c_�$ީ�ЯdL�޼;*���r��
TV�X��]��H�x���_vA�����|�
��>�Bo��Q�gc2��D��N�h:�?��ܳ۶@�t��B�_F�$pv�fۥ�����S�P�Qp����Ϣ�U8�Y��Dm(\�H�ʓ�^Au�?RZ4��'��cgl��_�W���!`a�+��U�'�1-��:�7��w����C]%_7��涻PDo+��sv����nF�͏�Cd�#v��&r'y��C�iƥ`�b6��7ٜ�z�\|�J��x��|�?�#�?��?
�&�=�
ْOa~9֫ND� 5����׹�yD;R�2��ā��t���Z�5<"m�Tmu;`�P��yT�6c4�֎p�B!�8��Ė��R�H��v��]d���K��k㍆S��9Ǫ2G*Ns�҈�U��f�|�����*Jr,@��sy�C}�d�W 5�w�A���h����?�;�#|�0�V�./1+�}z��u�ҡ5̟�D:�