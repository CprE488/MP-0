XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#�骅f��4�.�8�؃ �m���O�]�h�1um��1v�D׏Fz�м��jq���o���q���`��("�Js��R˾T#�T-OzN(�@r�TB���*ʟ(D!��W�_�ǜ[yK`ܼV�6}�|�w�S#�����0
yP#m�NQ�x�tV|T�	��خ� �"U'?%��^�a�ʨI��Ũ�0��ʡzr������v�fK�Y����h�:,(U(�����!�ND���l:?��֧��[ ��D,U�Q��SB��1U6Q�/���e��a���9hh��7�_8*����Ib~	��{$�&���/ڵ�Q#���@}|�MP+K�`*&Y��ͤ��<��f�)X��v�7_���$��tV�)������LW"�B���{�a��f�9�����Y�.�"�l(��]�[�jr�zE�lmV_�B�f���u�gr�J겐����DA�[ ���r��9��J�Kb�F�Ú:����ѩb��!����yp&]\� #���~2�U�[ꀙY�s��#���W�+��w�V�V�rͳŸ�+����4��ms��c��Wcu|��y��
�y��s���`�G���X��<i��ܩ	�*'�-w,&�s!R_cǖDf;���|�K�v�̼��(ј�����Ě|7:����I�Fi4,#�sE��T,f���D�ٴ�[x���+~"ܭz����rR�^��SvF�ѵ��c�,���������`�����0^mXlxVHYEB    3fdc    1160q��֝8W�tDjX���h�pƚ�`�k�&ٝ�T�m�\պE�t������?�T'�ˠ؉�}����)����8_f��Rܸ�I�%}N)����%��BVmH�N����%��!B�F*4E;:�3+��gCɝ�l��C�yU	jW�i�h6�J�w�QP)A�Q�b�.@:y��`��U���}�09�3L��>Rj=��=��ߋwੑ��R��*�j���`��8%�v31&������9����n���yD�%�%t*��ɴ��޻�7���O���ՠ!m&�K��������+�m�;UΨ�`D�w�N�C�YniX�i��ӈ�~��a�$�#d�Sq�cb�xP�_uHçF�ⳬ~�XT�#/�7�X��q�$8�t�V��	7_����+�q������n�	���n�!#M��$'���O&��J�Pj�g`�V�͈<n�����W/{Æ�^Nh��Ji?�K���v���!�߬2������)�'�^0�����G���l��ӹ��ގf�\��i��;�-�T=�J�ˎ`�d��B	��ᣎE��Dn���%����bM��T��iI�-���ee��������~�2
��v�Z�U�x1��n�����B���Ӫ�(��͘栍��8M�e>�b	�L���~9�ĸ����]�j�X��'��r��ּЖ:���+#Z�%�z��16��^mcR��n,b������Ѷќ�Jn����X�0�\��3�+A�V�'��v�c�e�F'H�M�λ������u�ʹV�5y�\X`1�	*]��V��֑�AV1|�!�����>��IKN��-��h�]b�F�H( P�}�h{�n�iL&|*t�.ݩ�n��De��djw�͔�s��q�Ϋ��珞+��1c�f���ᏻ/�0�L��n:�����rL���QN���!�j��Ǝ�����l(���ԡ`&�!�l־���L�
��7����Ak[n��i���1Xh�W�Y��$g���['�Z��izٱ�]o"���E��j'�*�:hmN��}I��tU�����J�?1c���Ս�vO6D�5�^�.�}���Kz_%M	���mB�	�0��{��������ְ�듀�ݹ|��9�'F�"�29�fi�6���x�+v6�a����s�'D6r�A9|�9�*3'�$�����ޗf�:v�<҈�[�L�����[l�~a�'�iD�J�ɐM��(��7���{Z�=푟�|�W^��`R�Ś��c�S#���#��8p(��p����Θ��&s�	S#�k�W�֬�=gf���	��:���G���wySZ!^h��K(1.����EQ����t�gt��������p�rX%����p��z��	]����s�-�Oǟ�wY^jT�;��E�nA@��&�V&�z ��W+}�����*�	�%A1Rd��F|W��W(�R�>�@��%��?i�C��^�K2c���>)g�����F�������@ J����L�����o�3@ݟٕ^�MK�S[�6��(=52:�e*)C{d+������ҋ��7��j�Z�E�
I����[h�~@�\�_�I���Ta��0A��	t,�4~�+����%��%��Wߛ�4s�H?.a�3�Ӆ��������}?A�P��{�J|�8��2y�s��[	9) ����_!0O [���3��Z�[��V�����'����bR�3V���?$���C?��偿g|e���ڿ���=]ߟ��C_d�#^�������wN�Ϭ��v<MQ��qQ󭽎>
ץ&�!�����!kJA�z[v����(4��	�/a�M�)���4,�������x�+�:��a�O'����{/�4�UU��jݼu��+��]w1��5��+]���c����,;�ew�9�R�K�Y��bn���<��`I'<����}4ܹ��U98'��Vg��gk�S������nm���kn��G=�Ʀ�o�R� #��Sb�;[l�\xQ�,B1�����7�|<�Ph�뼔�Bj�t���fdj�+I��4�T	ʁ
�!�$#N5���&?�c�w�=��Ԥ�/3�ZFŕȾ=)Y���C�9,�':�&�6oW�>B��9�5m!H�L�b�U�
0ҧ��r[��iI����5�'	��,O��%	��{M�f�FϜܹ��.��U�D�ql�UB���ͥO:=,�Znb�o�ȁ��R�\	,��]@�Zv���q8��Zl�2�cM#ۨUm�`��mfa=�Y �"���`���F{~�o��;4��3]pFm�%�Oh��#�V�Տ��Q����?�\��%Sl� 	��j�R(6~�Y�@��	-RuW��ݡ=�oSݗ�M:H�3�II���)�C��$�9v���@��9������.�#E�t� �啛���J?�vŻ�y�ՙ2W/�I�0���t��w�yp����7f�BX{a)U`������^�CU��|V~K>��8t��2����4���ڣ����O�%=��fL�yd�9£y�ۋ1{%�v:��K��ے��P+:�
�pEa�ʱ'�:_����Y�0o3(����NZzIb8׽�+�L�)9��k���Y#��f�V���9 ��Qp9��3��k�	��F�؃���-�m�PlԚ���(�^�����Fa�"]<�`�V|��`����Ԭa.�)������pt�����e���꤇P�l��I\ ԙ�^�W�f*~}�2���t�ƐqS������g��E�qh]V��0�������]~w�>�{>�q������
.�P�;�%�Sr"�n+|`1�ZtDz�#�x��TU��;t��(�v��+�Us�RM�ےta`G�g�?�7] ^/�X؞z��\�l�y�/d��ɡ��s�#a�����ؼ)ސk�Ѿ�¸����0`�/����,y��Ȑ9S����d�?m�`v"��c.B�Y'f�c����xKIJ~;�4���V$��M��W�as��з�'0h~1 R���o�ɱ]��e�����&��ĸ�8��A��IY��e��o��G��Ǵӿ6l����x����*�hQ�I��ù��?�YA��RP����b3�g��I>St�?��"����V�ɣV�?����1߻�s(�gߟ�*}���%�ԁ�T��+�=����O�AA��Re�E�p¨�Qhz t��#�02��t�
{���;��"���㏼�9�q���h隦��5W���S���\���#����xdM�,t��k�p��f"~�GJ��'P�����g�a	Є�2P��>�vG�'�7��4��جHwU�C.�G&�/�^��ۡ,c�����}7�s;X\�^r���a|K2���E=�!mc���S���x�S$��뎇Z�(6��������ؘ�z�'�U	OKTl�*ip��<#OWO��*��^���e&���� n`Q0�cZI�}��I�-���}D�~�2fb�rx��B��6t�יE�D�Į�o�>T���מּguf��.g8t<���'fI�MQ Eg��g+��P<�9-t�*������� *?_��E��3�e�9����؄�;����M[��7�]tI&�.Ga����M�CG*��8�6Z<�R:�m��f���,*!�f"����R"�I՟�P����E��֕��l�@���  ���@��T�R��l�^H-qH4hb��4r/��t��^��n�+�=�8,ª��Ō����L��4a>?�n�W�&z�����<��j�_t�ۿ�R�R*�5��	��l��T-A;7@�2�6w0�h���fm�}�T�y��Ի��C�ƚa#��0@�ʮ�~Ti1.�9��Sվ�8Cf���z�!X�������[�˒��j� �y���������h�r���J��
[�ve9kp�:��a���pʊJ���V?��[*U��	pxI��~T�$-��gC�ʏ5���e���R�zp,(�߽�C��D������)hm��7�3����w�RO��!���x�1D�8��}ʰ������m\&�5��3�V*�m��w�L����eS��PS�e��p�E���	�R�O�>��~N8I�	�Rh�;���"Ἔ=�N�̩�D�r��R�QWDU�C�v��Nl�7>^JIa��&v�EپĴ��G��z�}��ѭS��l�Sq��e�V�������H���S�4�{����eû�����F��|�o�C��,�_�R
.��DSQum�/"%6/���7:j�U�!����a��@�߬{�6\ �ѱbܓ���4�`r�w��mFe��M