XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���e=�RGE6�xI����&&y�%����IMR�$��m�=h�68�'�̫�ɞ.8�k�C�c��FqԼ���V`MB��/��':�������i�焮|K��e����ކO�+X�h������E�h�;�Jt�������M�Br (����_�@j��^n%}m�.UV��.�$�^*(GNi��-gTE�*K?�1����g`j��]AbNef�ҝG!����2-fģ��9c��4�|�~��"���X�1�-�'����j�JA܂*X��_����d[{�$<;,��	8���]S��>22S,=��]�<�����8��O+�\D���W�@Q R��F X���m�FV�����Et�,�n��h�^+��AX�&�:^8P;�R�^�J�o����͙o���hBl�M�܊����hl��{����B¹a�bH��ڢ��A�t��f8���zT#��>\�D���A;+E���>ϻЎ|�����٩&���ӯ���2E&����A�UC��Rh5��+E�4_��C�$���i#�]�}v��ˉZ�X-�(N슫�E����х=F+�X���XI5}�(QD)�fS�<�$��h���E¸�z��+Q�����ȗFEe8e�\~'�SQժ��;��(��@;Є�!p��C5�&��6�J��Zg��^U���d"��R���)5O��j�0��1��6�\t*�Ԉ�͎�IL8�}A��A��Y��Ed�q�I����XlxVHYEB    dd8f    2160�֎-����e�.PR����wMj���q���Z>����>���jTr�:� �*ʂ��N��K�C��](�����Z
�s�hx/�-�YQBK ���d��t�� H��:�/*�Q0ꤙ�p뤷n�J�*�0
��2�����R�U����No�����K�ڴ�Q�4��Bz�>���\�k*���0�_8 [����!Ӑ�dRS.�)Q)& �ThE�O��Va��/EѾHN"zY[���4-M}
g}�˄�s&���qt]�#aKWd�d��̭`I��oӎH)��晑V�\Iw�\�Hh�7�Nkb�,K��>n���oq�m�h��X@ 8[d���V!�V)��[da�8�Fy�t�'��T�ࢻ3f� [Fʰ��x��3�ۛos�h����)��[P��O�ȯ�i����m3,�n*�����j8�[�d5KS��<���D�x�-�8%�!`=��F�77?7.E��P
eL3�XP�a!�#�Q�*4�?�?��y����_��nj���D#>�V?% ���1И|���Zm.�?4V.�i9c�A�b�.�l��e1�mI@K�^|�|��QE��c�?�'��&�v�ֺ�=X���M�k��h�t�S���`l÷R���F%㍔W�^�㇋��ˎ�\N�v�VG��"����F,��uݯ��,�*����mXc���>q�/�Vu��@#�DϮ?>�߀�凫7/��UF1�B�����{%T-M���sx�bh��Qm��|̩H�^^ <��{1�Rf��:g���|<��ZR����n��l��m���s�����o�ʣY�|ef�O���.B�]�ax��p��(��.�X�I^��Z��zTlS���,�cAWٛM�j.`\��؆q-�x�*�n�hf�܈��mC�֓��w2sI�w�dP�@r��Y�s(>]Zq�I*yKoIm�bKR��kp}R+��	.�*Z�g�C�B�U��٠n���w\gkOJ����hP6��3H�s����X�p�П�%���(�H~XR_~���Ƒ� �;��V�`4��{--n|�<�˷�X@o��m�[�g�	銳��4^ŨPug�Hn����T�kl����,���������6i�>�y:�4�}���t�2w2�g��Q�5�-R �Po�ʇ�b��{��'P�}���onO 4D�9��\��Z��0��@�뒂(^c��,�s�9��Â9-<���0I�O1�]u���洤@e�����H�a=� �-�2���Q� w6}�1'���/�pA	H$��?�P��O��T�Ĺ ��
2��
`2�Wnc| u|kn���3��	�KCʒ2��՘��LB|��I�B�ođv��r���s��Й�&�l����p����u�![��꿳�lr�v9��|Y~Uf)b��埂��I��$+,�3Nl�����F�0�{f����Dcm�v��ȯ�LZ8�]_����z`���\!|��s�w"�[���#� ~��uQ�vq�K]�&��D� *�����L����Ŀ���#�
�$;O�p��i�Rvh��ݸ^�A''E#�*�g��q�N|s(��t����N�p��f
]Y���W����u�/U�^�`���	�/��/�H]L�i���pO3��e�z���:���t��,��FR)���Ni���>}���t��Ƽ��}���^LqrH����0�. �]y�(�Ta>����Ǘ�Nr-�K<�ru�K�B4�V��2���f�\���i"\�s��,ў�5&�ɃM�CP�}bS
�e�Q��L�}������K�Sp�7��ۑG@KA'o���&B�w[���P .H�Z��`���	?���� w�8���S�
���hr��!�Or(�z�>y���.t��oʹ
[�,�,T����4�6��n�hNlPx�%)�9�/��o��0@?�~/r���Ҿ�T��U�m$�B�a� Æ�7�*ːcG���(<�ͨ�㝚����jݽ��hX�wEm 춺�v�SѰ��޼���k�K<q;&4�6'?h�Tod�W��_y����1O���c�6��sqY�������46�ޒN�&k���Qc]�N��d�ʻ)�y�:a�������H��}�j�ZOB-DEk�(X?�����a�A�F��If̖��p�oAS=�ѿ{G���CQ��>8�d���cYc(��N�?��үd�TZh��5<�z���&�.�5V�7;���3�1��ִ�(a��A���$u����6�����q�>)��zv�I=�4����^Z�*�l�n��+�"ˤ�L�C6}z���:� G���ZAF�x�80�E������t�~�A�Sɖ:kx��x���\L�
�`��2K��T�)Q,0����٣�H2�;@>���X����x��+����ȴ�J�C]_���붸�ٹ&�Aa��l�J�"M��Hс뙆�*&��|"�hmi_�\0�P��K�|[�	�7~��O�� 5�3�.Zf#SS����Ǔw����kl�P�"������Э�@*�,͌|�����6�T���?����?��Xmk���?Dѻ3Q�Y�L���./(|jeƹ7ǥ�s��4�.i�ҹ@Q�L���0�v���`C���1�/\��ly^��3?/�]v�)_�z{C/K�u�W�z�Q3+ ��>�?Q>:{�C���%�EZ��$+�Va+3�7�ç�OP�Uε�Rtj���+e�=#�l��"�����p��=��������{X��z���x�㸩�Jtk����J��s�Ѳ����%� �x�8����{�b��[K�
�V���+��S��+�XL����ú2@�p�C���h:�
#���]wd#ڬ�}��$=���u����f�w2�Ť4M��=� �Cwj��Kg\��It���A� oӏ����}j�Qq�Q$s���D���ɾI� -�����5ؘh�{�e��%������K�B�Btn�Rq�"�<ɢN�鴎1�z/����\3�m���b�x�Qro��9r�c�2� ��*��à��s��B���kU*�ؼ��%�2�*�0���y�X|���i��m�8�uL`5�moL�v3wn����\O������tKh�����;�>�
�RB�XԌ9�]��f�F}��X�_�ҎJ�a�{;�*!�R�R�~�����U�X���gO�FүZv�f���2g�-�k:��8�粵�v�;B�'��px�+��nՔ솦[	 ]u�	H~�`���D���VK[�֠Ԭ;r���[�(�H[S�S��?C�3���ki.>��˲�9�}"�#��i�E�2_�l+�֝��ϴs�iH�joY���8��<�y؁H&2���+\�A��,s�k�T���s$�ڣs��RZ����r2zFx�h���{J1�y�D\`d����u,,��Y�m-����X��A��On{y%b/�(��i{����Q��od����9�*���a�ye�/��ؖ�Nl2�W��,�{/�+0��VD�F7ơ�a���ą4z�]u��"���T5�+ߨ�<-���u��(�tv��_x;2C-��r��$\ݵ]2�Y���߁^?�eL�"O���8�ewX���h�.Q�.˞�oq�:�v4!p{�E�ߪU�:���A-o�R�P�i�Z�I���I��fVq��Qǋ��?m�[F�U��m��!Wx�Y3�8Y��Fe�K��I������<^r�� Ĕ�4�=Ɠ� H�{ڹ��~ ��=χ�W�B�-��U��țE頁Ӥ��?�C��"i<oc����w,gjQ�	��2i� m}������)ѽA����Yi�]*"L���l��'�)�9�/����xL���6Z�X��� oIA����!ڭ�pFg�jU��"��XY!�ԫ1P��gl
Ϳ�;B~H��+�}!�Z�� �Э����&��jK�1 /U��e߲9�|g�ڞ�k�;lw���#R��-�)ޅ]���?�מ[;v�@/�h	��1MO)q����

R&n�/>�M8��L�-��ew�L	@ZH30�3������{���O�n,����R���s{n��m1�e�P�q��T瓛5Er��C�k��U�X��(Q1�.F0�$'��Y�v)�3��{�ۢ*�=ER���N(a��M��&�>W�r`�	�p_ ��/��[>$r�Y��YgV�D�/��y/��,��Q�Z4n��)[�*-_�D�Ņ�H(J�h��<؟N"+IL��].np\Gؐ�a#I;xہX!�xk�O�=�r�m��J��f�xG޿����'�в^��ߘ��E�Gޮ� E����/�
uz
ex?O����`5}Ԗ[�XG���A��!4)|�fHE�� Ǫ�)��/�Ĉ�5Yo$m>A=��8�!��/ì��r�;�Y��P���eTw-��>��?�����#���.�gDanC>��_�IC�I�'�U�=����'��|��O�^�4����
��Y�x̰��b	��{w 29{�re��T4�g-�����/]�[�R�s��82��9�}�}��μ���q����yJ�s[���,��O3/(JfJ���㓻�:��Cx�b��3�?W�4�J:����ׂ�e��/ ?80ȩX�(�e���7J�)!��q )���&��(�;������P�������4a.�t��}Xk"��u8��\����9-ҀX�N

Tx �8��[߈1OV�9=}@���d�N��9}Ë纰9%�Z��`�W젖�qX0fl�U�تo����� �b@���_K�j�
��$��a2��������8���BW>�U�D+m��x����.�[��^�"�w��l��0�ȫ�����VҸ���3��>|�� ����0�؛�A\Lx�,������}���l��H�չ�E���=$6�X��-��0���5Ylv�ѓ�>E�;�S6�;�	������8rL��^w�F�P�o�v�ۗfn���0���:�{FE ��1���Wb;٠���k��<��zyt��&�6痙PU-�0���o�?i4�u�x�j[]�	�������C/�����@W�r������߂���E���ǂ�H�~+_���9��x��_��E*� �~�}��8Z�AAr.Zdڐ���B��!����01���iN�W��2)�=b��y V����<��H��(�V�;���?a��!'���
�c�|��wE�E,ߕ�엵�E����z�v��!��{+���xA�X ��p��zۺ,���͜�#qdqu"�.����G�,	T�g^�i��m7������	N���RUi�
��H�Ԣ��yĔ
�rS���6�6�6�[փ߈�m�yZ��g]����1�or�����kh�་!��c�����=�`�E�ia��'��Y�neR�i<�"a�93������Ӥg/{�Z�@�`F�t8���ղ�V$u%NG5=ݥtY��s]m�_�V��V�p��,�}���*����̖@q���x`JW0���X��l(ye�"�A�mQ�2YSF�|���YZc� ��2p7�K�1����,X����}�|�Ǟ@b�cu�{�j�%`��s��g]_�B=�.o�^�T�lĨ����0�U+�j�2Ú)梧
����0�I��+0�ؙ���3ޜ�H�ֱ)x�Ŀ�N:��$<IlAGs��]�g\�@D�`���/{&Q�[���3�PM
�u��'0A�Ūd^{�Q�����l��"7�n��J�����?Y�����^����l".�0���5�/J}�m%�R}�%���D6D��͍���	p��o�i��'��5�YLA�>����V�R%��7����~s�L�N��/�� H�vŮ\�v�<Fu��T)�VJ5 ��xm�*��m�`��8�)Z��Rмl#j,[���Z[���AT���$Z+����'�%\�^E��6&�$��#��~b��&AM�C��{��z�{�J�Ѓ�)�Տѓw�e��s����R�<+�E�@O�	�sF"m�_�^JY�':�"W*��b���@@��(~�r�&x�]��b}f��of*-�HV��B'����Ș[����N-N���jq����F$���I}�L��:KV�$�HI�HBEU�6��]�(� '={#���bAwJ?[����?���Ȥp(� $$uMhCR7�Ľp��zkky�G�m�'�{�3�G���W�{�Ţ�x�#f��ٳu�E���q�؟����U'��w ���ϭ�ى�����c����0=�ح�������h�iԦ��e8,�[)K�n��ʏ�`���ht�M搽���W��5G^@8�c ݤ�H2���;K=�v��fJ�'OI�8	o�wa�S�+q��8�;���}#u8!��DC��K��rR���a��$]��Y^�'G��H?[5���]a��C�v�}3��U�N�;Y��C̀����e��-�~�pP�D��1�[��k�|U�f�X��B��pM��0T�{��� ���N���ڊ����5�!����?���F��5H�?66��/���%!��&��ARJF5�]HXX�m�B�lWBpڶh�䆜��? �I����������x���"�!dV�^�K�+�W�1�p4X2�k�&��nn��[Ȗɿ���N�a�IН�)&%h��!6]��+o���h1庩Uif��~o�������)F�X�b����9��F�����]a�[����z�����n¬����"��M�ٞǒ3}�C�N#óC���ĸ����@��1B�EO�,��!����9�L��O��V�Ρ%��5�	S��<���L��D��賕�%�q�=y�U�M-��?�\�A�7����@F79`^K+��۞&<oz�������x��A$�`a�ޑl�6����Y�,��48I dvl�ډ�s�O�{}��K��>�j���1=��,��'ń����\L���j��� ���eBţ}�F�ۥڠBW!�V���n�3�d;��_Qmq\c1�Q�s�р�81�.M��E��<�A���c�ww|�G�1�B3Wg������*0��9��FF�N;��R=�0��ME;v!o��&ҽ��ùIB��_�F/�}Ɗ�c�R��d/��y�c�'��P�<AV��bw5�j	�5 }1�"�Y�}i�<��B�;n
���d�q)�D�>�D��Y�Ϧ=��֫y0N��&���N�n��	1ym���+J䈅I��? �SI��2e)V��zx�#��VޔL���|B���Q���
s�'C�+�h�͉z�� P�����+[`�x^%��q�j�,Cџ��:��'F��s�sq�t\�~ܳ�:��C0��ߠ�Q���+��	���$���s?�e��o9�����[N���`��v�t7����h��B�I,SV�"��ۿ!�p�*�eĔF�r�Fx�a�-_��w٣e=�Ϻ�LpjA��_��HI|f�rt2^M�Un_�hI�qYFʢ��[F蔵��=~�\SCJe�-?�?	�0t��K׻�[����E�jQ�|��(Z^|\���6S�������i��8���m�y��!u�� �+�o��km���q��d���j�:cNp��� %��(?��x�)FW|�z��w�wć��&ڋ`s:To�b��N��5��/�_!�Jmӷ+y�T/Y	J�����˹�ᵏ�.�)<3�ʘ��/S�q�>�,)Y7W�~�I��5�:B�[oGC)L������=�=}�[��نd/|��Wg��Y;պ-v�Y����: 4�p}52@���	k	�s�ZMH�y�zuL����Dۥt�ǟ���*�g�'�Z�A�w��|][�xz�2u$����nGX����҃��A]��7~�֚��ϟ��P!� ��m6��S�X�Ru�W5<�E�V�k��|V�/|���gƏ�c��'8JT�ύ��sɈ�W���q;ᖤrK.��(������L �x��ѧ���B��\P���A%o�����
N|�ᶱЯ��Њ�/��ǌMDr�;-��w�Pv�	7I�N^��<. �P!w�j2S�$Dd�v���_�BT�*6p�W-���M���3���!���F�],�}�ȩL�"5y��`;!��6����WQ�^�Ǜ}f�"�~ �16��S�-NFƤ:�z6��U�p��!a�׫��d��ygs�o��
@��I_]]Lf᚝@�<Բ7_�:�K+��*O�W��1��n71����\����.ի�W\��`e�i�L��Ư�T�L��J�ɸX��>�IW�Ȩ���Cd�J!u@t�U��7�W?�+-:�}���C����<
o߆&J