XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���%���܏�%��6w9V�q���l͝$R��2P[R�f�o�i��%��z	!�s�A��t]8B*Gx�����"VSD�J��,ۍ�z�y���(�S�����,�����D<�2G�K�ZZTg����&27�qӊ�p^�؊V��4?�k ��m�+�]7��z�Ҏ�)�@2OY��;"W	����R��zP�rN��}�v2���#+��
�e��������&Nf�o*��/�-Ӹ[����k�o�h������s
��_
@M��w �hG�{�N��CI���j��c�V��3lh�b�-�N�N�av�,��":#��̴�J�|�3��X���/]�ǯw�P
�����(!�*'�����Fc�����Hc��s^F����?���� ������T��G���%���3��S��>���D&���`����cv	�~��7 ~�]fO�$>�˘G�C��L�a�^ǴL;Ǉ+@R,�z>���{ɫ+jP/�n�.� ,M=+ ����E�����v�8��T��yY_�а��7Q>���!��S��P�<I�fz��Bm'��6�"�bq�#���V̹{K]�SCz�4�2�K<^�؝)�����6r�)�! �լ�_�Yx���v�g�:#Xx�p��2�[L�<E)B��c�$@�c�o����������h��-�`��hɪuEǄ%J��T���l�j�Nd3���.=eJյ���љ;��P�F�}�XlxVHYEB    6346    1790�>
�Ahw���^��aC�����fST��������H �RZb�G��z��V�~�'���j� V���K5�S�(u�) @ ��5gB5?�]�kO���|wF��ƣf��&����-3$q ��2���ކ�i���B=��cBO]�O��Ս0��I�0D�3V9����;�ޅ*�J����p���e\O�┲���h�0r5����^Ո��f�w��7��?�Z �G�׋�-b���i篏S/���P�l �Uٞ?�ڰ��I9��[2dq��5�+3*ȻI�Y�.����`?�2�8R��n'3߹�- ݂��mX%P�p�}�.��2��N��Ln�OM2|-�C�����So֥�J0%F]L�59x�H�>�ҋɧ��-(�|i�g&�/���毲���8����k%6	���<�������H#��񑞒��Iܸ�U���T��"����쏘kM�'-3��1��5�΂���y���c�q�D���t���9� \&��Y�H�T����}w�8�|/Yq �J�b�INm�w?Z�ڷ��ν[l���NzS���F|���Ј|'�o�0ޤ��:
Z��<E�Z�|�Հc?�ѡm��]헉)�|��C��cܾ������U6^Z.x}�_���$������H@�撂(8#5��\��#�(FyE���Q['F�,���?�|�0���*A�*��.^#L�8IG��C�Hw�̊:׾��~sw���m��H�[>g,=x��r=r�Y�>'[�%��Wv��7m)Wq�����o���&�t"2(�6l�Y��G�ê�$a�}�^I���4Mq��)̰7m��KL��`�	 �4{�N���/������u�'Z��L�q���G�e�PN�|��^p�Uq�S��=���3`�x"0�إ�������YL�9�~�˜�����ڣ��f2���ç�B��A����p�m���)|8.�n��􎙎���3��Dfx�|�%%�'������&/�؅��n[;�*gd$�W�1���g�D���_�<��g�i;C�=+�o���?o���F�YG(#[6�����)q��N�8}���6ӪŰ&l�.R��%Α �s��F���Ņͯ�j��qk�N�t�g�"*�!gu��Rvl����i��d��ׁ�?Y�����9�����ۣY�����u��<D���κ�8�(Z?� ���+A���
�hG�+l�`�q>Ǳb�<:�3Z����ֵ.�f����Z�
�\�m>c���s� �Z�
C�*.�_Φ~&w"M���c�I`IThkQ��p�c� ��a�{�\=�*���ɷ���5	4P<�ʳ��.��h��e�T��M��{��ز��>���@¾4u�1��ڞ9��W����!��-2n���n���.����O�����{!ʑ��L]�V)��eH"K�I�sv�|��k�?$<��>o�~��{RP���f�ik郁q|đ:WD�*mm���)ޖ�o��L+UƧ`�(c)�TV[za��W��� �qn.w�$!+�/d��$�~�f��6}j9v9�,7t�V�ֆ����/�g�{��qq�f ��{	���Q0��'}4s֭�S�~%��l� �U�a�al5ZhS̘ �;1b��s{�<�6���GE��ڣ�K�p�a�*��}���ڏ�<�&���X���y�Bx�̢�o
���(���!Dt��h�l���ke���Q�?^��-��u�C��3��w�	��e�/���e��zzL"_y�e0��tvI�̲�V���.7(�W]-��}W���o��܊�0��1n���s�OAi,�7yNC�,C�5���)�E(�6�I���)K����ε�k�
�lNCcq5E�p�È�~��h�&�I�e��L�[�cE�ՏK�f�O��/��a�hc cҹ�"�ý;Pǐr�<D�p�J�z_ι��P���m�r~^t׏*U"u�
6ie�?*2�^k�83��P�i��s�e��h㼔:� &^��P7�)�,FnQ�Q�f��깫�97�rR��%�<�9�0�׿��
w,��d@��8m��<Ǒ�&�w)�wy6�ŋ����5���Hb�z�C{�Š8����ۊ���y�a������0����n�ՙn�[���+�$ރ�z�~�-�>1}4!G��:��th;��
F���G���!b�j��P��۾h�W�c(<j�i��/��:�
kmv�Lv��`�xqI�U%2j�|�$=4�_��}�{l�ہ�V� [ѸMT����%���C���}�t��)�\4[��BH��T���g��Z&�3�y�Ne[!-[T5���'P�����>�O_o�9no�����oZэu�bߒBw�g�I����
��1�i�I�y��:�����`'QpX,�ZWЅǚ�U��#��=�A�Z�b���U�qa��Yj�!�X5���n�e��u"�QZ��x
�?�ڬ�a���?��<q�H����QR�3��SQ�#�з��" y�FꑸF�����<_��4j��t�rzI�\�=P�.?^fQ�m;�jO���Iu�����<Q6v@Ŕ�}��(�'����3�n�{���bLS]4���H��I��:���G�"�`���K6�$_),H��јe �Vo�؟��FAXz�0 ڒ^ (���:�F����֌�;<,`�V3h<��ARk(�!q m!��%��nd�`-�8Go^���۽*��̲]��W�`��y 5���7\v��Z?/+��3TU�~hx�F<(��"4�	5kZ��wN8��.~m���&�Q�]��}�.�dʷ:�^�^�qTdW#e�~k����u�$�~�J��n^��K8@����˾�AM��xh�d_4wY�e0ѶI��ƗF+����2S�c|\l���֪�CzF�ͥ�to�:o�ߚ�����ڼ�NC`�#"*��5��'�癐$���g�+�0��>PO�+�{����+h�-:�0&�Uc�Ns�N��8��-���_��(��p�#��"��d��N\����fF�F ���%D��q/��b�au[��	��/�ۡU
Wg��F�a^��:�>�\#�U}���]%���m\�-Ʉ���䌒��laMS���>G���YK.1��(��lم�<_�s��"��Ei���;v�NeFP�Q�X�9�M��{�7Og�$�OFݕȐ\w�q1`��B���J�a�,6H��w^�u5�V�@N�ͣM��!��l��o�1����?�M�z�k�7*�֤���zu��:_VnYFP%��<m-�:hj�O%N�����؃�����P�U��?� �
��*��N����=�	1J,�k�����gr��_�I�k�L9�:�(x����6?��BI��m��g�p'�
��6B��KYؿ�ڏ����eoՊ}�������0��n�������� ���	��B)v��g�ϴ�{f�W0X��B
I�x�Tq�v+��)l�2x�&� ��B@/�6������ΞF��k�JU$�|�;�W+�r��എvG:+��ޤ$���_�*�{X5e���#���%\�5 �U���Rv�WԐ��O�s�U���f��@��@��mř�R q�282U�Ƽ"�$���{Mի�nSsuT��6͉��}�y_DfAy<U����U���0-�W�.��k^�F_�2�Y`%��@�.Gp��%�O3j$��4�7)��u�UVbv#��+<h�L. ��������vc�.���@UW<�9�<݄��>qE�c�ƾ��bflً�Ŝ��'IR�I_����K�L���?h}�������#F^X�4Vv�)a��~ip�e�o�/�4kV--7�J,���5R���j��x��T̹��?��Y�)��N3oR^�nK%1Q^��|Q�P�{<��xF�Ad5��~ƒ8֛e�F��(���]Vc@�����K�<#!6���&���o�(Ekͭ����8�1�,��<�Lo�]R�ic06>4��������fU��������f��n��2����J����Q]�&'^�ņ[8����:O&�&D:m��l ����*������YJE�����%�g�/1FE�H:�'[�X�(�ӊϫ����q��y��٭qȏk�b��b&����+�=h�d��F��xb��z�VN+��'�C���I>{㢩T�}H�Q4Ā�>�J�)�0��S⦥O�F�* ��V*-fGh�w�����O�VS��Gf�4(-%���j�;֫�O	���.v[��0��N��;$���*>ҳ���|O��-/i�|�����S����H�L��C����T�^x�Izզ���Z��,����te��ʻ��-�k0/����xU���q"����)�п`����%��xe���Tyh�'�e�)��2����YrHt����p Ӫ��(*�c젤���e&��m��w\<\�YYp�*@(R[��G�am^fb*����d���M~�SuO�9B��]V����J�^���
��HwOM�ӹ\� *�QX� 'w!o��0��HXO�󒍵�5KѲ}��ݼ�!�&aS%Ua��ڕ�=Y�i��$||�?L��}fG̉�e�u���$,����7Bd�M��cf����!��z'N�\$��мոk�MٛwI���|�y`�[::���L%���ԧ	�R�u�D�6��C���#"#}㗼�D��fD���A~O,�`$Ǐr��O�r��D���"`�����b?y(�6d�8���Q_�]�����
������g)�7��Y�粼m( &&ړ��Ar�_��dcm
���]M�w�=��Ӧ!�=��3��T�I�u��=�pYL9��qR/���h��1���z،�_������xy�:f�,�mNK�~LD5-����4'u-��	���ΑI'�!�!�~O�&?�7ơQ�N����n3���Y��"M_��7E�L�G ]:�+z�9ۺOl,�^i{���n�VHqw+1c�F��׌}yכ�	!]A����l_��(��V�*��u�������f�Ά��B�3�I'�'�ge��Hs��S��'qQ���V�y� ���W��r�©Q<���D%�#��V�/��@��!f׍O�(T�|Je�Y�{s���@��J�h ������paE�n�����~����7K����j�%{�
�Y��ݓ�uu�:	P>Mg��`�tO�-4{�x�E�H���e�	�������y�S�)k�3V�G�9�����q���!�)z�o4W.6���WzXi��<��}��Wk�1�����'O��X,fUCjΆi_T�B,�J��W�v'P�C�A���&��

4|�IØ��!�B`���',���'��hC��
Կ�
)x�S�8��
g�C��[���a�����O�e���h��L�[1yr�5��m���j���l,�4��3�>��p���t�K��=>��3���ɼ���b����̻M��͵�U0�[���������s�Nf8�ޟbl��4��E|�\lF�TIL)�Ìr&S�N{vD!��j�������x�Tɵ��w�<�]h�H�Q�ð�AE�(N�ʵ��{�K��S�P��6����gD��:� n1M�\z4M�]=�E7D�`O�U�����k5��Fr6�6?�A���JC$��i��lw!|��̠�B[?�S�#&";�9ۓ M����4�0���e�@␉tF{�.q�.��a:� *ԭLߑ�h�X���L�Y�Ɏ���g0�Z��1Ȝʋ<a�?�="B댬�=$UȞDt�S)�Xa� �˾/�E�ru�oس H�"A�g����Fj]�φ�H������O��Md�^�3Ř��)f'�=SI���Wjb���оq�2�F.6%���
��ɨ�*��pF �3{��}e