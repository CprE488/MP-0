XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��s�U�5p ��v�;UԎ�Tb�����t� �7�.�v�]���A�}MGs�ff�����;���KH��Xsx��͋,����D"�k?^�}��S5�lU
="h\U��^p	��[�a��7ຠ�Y�Le�Ep�@�a6ڐ;��R�/��{�/<SC��`�=B��K����i�h.~��"��(tE����BӾ���o�{��\6�D�nl�
\9;�$�� �!�5�
�ha dp%
1��=K�DR���E�(�	�o���e�}���P����J���
����0K,��o=�)9�d��ة����Um�MZ�u`Jjuφ�ᨶ�3g���c*u>�q�Mn� Ϟ�;W"�=?1,��6jy�Y��'ŀt��:]����y�vzy�9B���O��H�]H�c����N<p��*�^p�������R]!��'b=� -����/ު�MZ���-�e�.��ׅ#MZ�
=/�{k�&�m��x�#�
�<e�E��
��f��֫1~�ݗC],�hۻ��4ي���D���/�_䈞�[Nԍ��1�����{1��s&�0wr�;��ɳF3�f�;Ўg�aLV�Kd��^�Ȗ(��b9�����g����\�	Sৌ�Xl�D\ȿ���i�e9��<�AS���.�w���i7����Į�.��.��B'�C�*��\��I��b�h��z�`�3`b�&�)(���⳰l���|S,Q����sT�:tƏ�d��큣 N�糨-��XlxVHYEB    42ae    1110L�?"�����L9B:41%w�G{NF�^*�1�.8�-�o�s%-Gf-I�a��f�J8�p&�a�BwId~���h�����(������Ā��-^$����-4���gc̀�"����&�ڏk(�RȒK�i<d�������ߑ�3誰�۞�~���`�䃐��a>�?�~�I"T�dgŉ���<��w���?��Aҷ�H�����}K���0����βJ�1�$��+3�W)vqѧ(�������(gε�v�X0������gz�&���-�e�Rz�((Sc+b��ڬ2�;�yN���w��㦴?�AMSv��U6CS�җ,����6[�̲�Y w��hݘ������/c��������.����N#Mj�ޟj�/����;�82��6X�]2W ��i<�u5��A<>kh]8���{�J'��G�Z�4� �(�X�=���MU���B.P�R�e�ڊ.�w'�[�b1lŚ�S���r����ӆ~?~m�K#bΕGO�~~�j7�����4L������/u3=2�Q�e\��<���jO���[��C�������uUU0-$�}l8�\���t�`�S�~*L��V�ͯw�3�2l�g<�.��/�]y�@:+��^��&V�MeXs�����&-����Ru������$�]�0���io�muN������3��Âq@�c��b@i� @��Y�=/�����IkG�Ʃ3�)�Y� 	��0�:z�r���Uf�:�[�&j� ��<!�Q�ş�G�0���O��S�1�:u�qw���>x������&y�k�FϚ������V$ &0���Ta�y�W	�8hi�/��'��_Ts�5hRb>���f��mM>�܁kqo�D�X��������l�f�6�+v?7[K��5�fo�����/f�S!���q1Q�l�h7:Lu�k���|'Ԫw=a~��-l�L�^F-��SY��U�'c~KvF)&� za�g@ή���x�\�t�TfA�: �U�����j-ޞn ����+��Ntr;�e�ʥ�U��f��\[[;Ԉ������X-ʷ]Di	��5�3��Ꮆ	3��j1d5��ʍ��M|�]��Se���������ۤa���#�i	�.T�qزd N$l~�ýM�De�Zt���(��8��4��7ᔂ�F*o�x�[�(�JH�lhƤa�Q��ka	�|E�|%�/{�6�Յê��	�{���䫷�N�Y+�u}(�!3�ν�����{m`��H�HÜ���KO�ޙY,��@�OQ��4�_������J�#�BuO��5�Q[9����n1�r[ @V�R�߄f0Χ��v���ɳ�%��N�CXt nA���2��u1J���>ϋ� ͜	4����l�gP��1����j{�tA���˰���
�f"��߰�~F��S�%���tV���S���q{/�9b�K ���)�bfL�Vb)�W��������'\<`��{ؓL���H�U�sMb����#K�X���ZI��z��-�R�_����RxE5�q�U�m6�n�5��0P^�e2��>Ie�P�'��q�]O̶Ёd1'��*!y�<]���V�^FC9�H�_�l{��:�ӎ �L�Ty��%��Ǭ35t=�.(����Mʋ.���VP����#�x-�aED���C^Lq�c�n�7E����=��4�S�:�P���6�[�����q�4�����W�,�g�SWPm[��Cں]�0�o�ɶ5'�,1ao= Ƶp�Z�Ք�O��Z2�l��� �;w�)�<�T�P�u�^"\�b]�~_RYxR�V싡�6���
b3K�)
Eʬpv�M@me�����q:�nCMz̀�n�DC	��G|[`�������Ks�W᩟jp�
�])]O$���H�D�W,=�#X�j8Q^fS ^�'�2��6�PL)0-؁�W7)�8����jd�Gᗌ2]�񛣀V�Rv7!F��|9���R�o �V`�F�H+C<��Rh,�����&���
�����+'=5�����9� _)�+�(��W���%S�RD���9ީ[z��wG�R,�0�{��*�M�%�z�+(^[z���+F�F$�@��ܝ�P\H����(v��;���GkW4t�7-�-e�~�]w�[�q�׾ib�睔�s41�q$�_�`f���S�"��|���="F)���樄m��\:��$z��u��rTd���@,��	+R|<��.�NU7?�Nq#�ڝ��=���6W�E�y�W�����`��3�Jxm�v�9_;�&)�t�eNk#�vJR�	I�qY��M���Z�Vk��6�|�8 {>��4�#�n��(��8-�����?�x���6	�ɳ�.|�6/�71�*lyĭ�^]�I,��6������(9���fv��ps͡c'���f��T����M��~;p���hp�\|�OUV~	��?��d!_O>'�L[(�(<��"+��Y���= ]�\H|��(hy�Űj��9�[�덁_z��7\�$��I�+����8EB��^b!����(m�}XѶ�b0��s��YJ�c����}��LJ»���<��������JYn-�$� �+N��b��G���ͱG�jn�6��8u4ƌ.�5X�T'T M�%!�����jv���I��s�8���.�U�������`��D�ٳ��6�.�E�*W����?������`��<�d�-����
�W�Z?E������	�g�
��l���p��s�Hg��3���y'��qM����s�(��U	�y��xX<���\�Ô��vO5��Q�耩�9q�������CdW���"f�[K/��������`V�{�$	��ڞJ�s�nn����%iӾ9�J��#0a�����w
�*�<wWz���{5���p^wcp(Y�����=�:�9�Hڏ�V�lH2/l<���Yh.W���'�^���l�(X�����a����L�:���ۣ��=��4=v�\"��\���Ie;�����Ի�3v/ť��5*5x.W�y��Y� �k�Q��*7{�*,�H��������l�����ӓj��21$Q��`ߢ�d7Yꓮ ����0�2�K]pVdᦿ{��� $��A����vS��2�v�$�4P�\�Zٱ��rA���`xΉ<�#z��ɗg��ן����
��ׅ�Ǡ�樑�U��z�c�����s	O���m���'R�i�"8���}�zc�K��ܝ�+-�=�}��I�G�M�J�Úg.ON�k|����c��2��n_^�E)gP�Q��D;Ĉ����8�	��ri�+�;5�-au<���1GҚ�i>B����őΐ�P��p؊�,� 5�S?��Xr�a�B?+mU����������i�yꌚ�?rK2�t��A��G����]�	a��$��b��J�*�g�RC�t���@��gg`��b�2z��J3�F�p��_mh$��S�H�U�8KJ�D��A�����E�o�bRH#s�_��c7�G>&ɚ����d#:9���X�2sg�~du�wDP�%O�T��SԾ�/���pm"���q�<�3Í���cYw�x,A`���5c���+׉&�+Gx0z�$+�'��|NŜ��H�ǝ;;��Y��|�B� o�(��Fc�`��u��<�*b�Ό�Ďp΍�%��b��N�[ 3jw�.T�L���L ,v����%`�l]!>��m�@�b�L��8�C8�ZfM���|�?�����B[����~^��Y�(��(,&�[�XTi�.$��:KhO�;N���z����(���"�A����x�<ވ�$�P�ݲQ�iz�L�g����Q�)��FU3�]HN�o�s�~ n�$ �1�:q���N,�膔�Ay�������
�:�א�[
�:�d�W]�9\M��}��n�/G�V^�&��{;���&�PFD9�_�3�ץ�|���6i ���F.%4��)�Sk���N��J�T5H�/�@��7�����p���^9Đ.��.�n�R�3�
�G}�FL��E��G�d'�輛'"��@��лy�9~�E�E�v,G����x�"Ҭa�W�h�}2�GF}��������+�FT!�u0�����U���g�=��T�,wT���|��Z��X�Kk�n+�w�6����J�Q�����0y�k?
SJx�z1@���{�C��
���ȅ44�����3��QH��V̽�o�����͛y�O�Otj�yG�a����hH����9�Q�Y�:��