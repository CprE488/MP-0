XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>z���&r����B�8�p���BE��sL�L��%Щ���EuJ�)Z�ɣ��͡K�4�\?�h/d�M����Hr�Lv���� #�^V�h��� m�����U9˼���e�K��1	����E���sR�U�tz6���! �2kɧ�rNM�EnT;��@�s������w�p�����e�Q�}#2iMv)�v&��Q����Yil��%`����2�\ 3��-�T^E�xL������۳�����F�wƥ��S��j�E�˨%��H��.�n��s�z��u��4�t�k��Ӂ�[�T}�U��	��������x��<�(;w�꿢�A,K�n���	j~>�\z������nm��?����Yg6�+�|Q�̻X�������s[T���T��A(~X{_\hi�6�Fi���w&�Pr�y�7�	7�щ��.=��N��z�y7���歵�$g��ep�m<��s��#i���$�[���-��Oȯ5^����5�(u�B��
���<��tb�"x�,,��X�e�ޛ��`q#B�¶CR�^�^�3�2T{P��̦qc�L̢!2�-�Jc������`��[â(�̹/q�*�ZzѣS��N�5�H>�u��4�4e�L�c��\nb�H6r����[�5|�&��a�M�"}\�`c��kKô���d�����O>ytqi��XM��[ܛ�#�k�I�wb�A�R�x �|e���'ጲ$9s_f�O���E�p��Z�����6n�(XlxVHYEB    dd8f    2160�:��:��HaP��=�se�f*~Fc�Y���[�]u�^����53�Z�-�G���m$�ia2�'���	�	ȉ��2�>���]�#qz���8�S�m~������棎�U��]1hW���f�m!"���n������#�ݥ���W"�6^�S�5���`·P@%��p;#1� #��5��Lk��/.�j�~$�0��GÚ�ʪ��_���=�=w�nr�Gr5ct	I2%��s3��%���s���^KfOc!��1���[����,4n�W����;*Fl���N;��^Y؇QY��Q�i���U�D�˅����svI8l}uj��㬆�6�Ms�M^�GP��gАa�����>��\,G-�.��M_�/��r�}�@��Ќ�*fB!�y Wn�{6;�c���\�1�m�γK5q����L�Y�ӄ��c���Aa�9�<a��7�p���W9�t�
�!eu�p"�d!#G��"���^'C��o,��|j����I�U�iWb����S�����Ŭ���i	~
}��o4�P���>���ú��xu'�do'�,!��8��NJ��ǭhZT+��MK1�`x�mUg"O����Q��T&x+��K���{M��B�"W�C����
�N}PW��R��m~������Ƌ�ү��>���σ���ʦT6�U�"�ϔp�Tu�+aP�zY� .�� �ɜ�������h���9�sJ�
"nm?O�dG�y�*}t���0���|��i����p�y�ZW��]`���w5?TGS�`�R��"!i���gw��z�r��C.i���)sXbl��w؋Ka��ߜ	��� }/�*Ce"j:G?ZA{�0{���f1�[~���fP�8�ju��.��3�Q.��+,j��*�����c�q��\K�}�r�z`\��? ��4�/�hy>䜯cb�Ƴ�>d���	���y��F�aP���s3�~=�C�GdU��`������[Om��v���q�4��¶�"�~��7Y��(N��c�_��]���:;��<r�`_�xDEGQ9M-�e�K�ے�9�㊳UT#mw��Z�X�#��8ÍqZ)��f�aZ��&� 5�,�//ȥkv�I_�%�zq��ݵ|�1l����IŁ"U|"�������3�'�Kڇ=H��Jv�g,�Q�W}UA����0��xfiksW�����.���}�홉��6�2@���+$)b��R���r��4��4����r�?���dJ�`o��Ib��Fe�7y���2�\.�4�Ҏ��*��u��(��OL�Z1�'� A͹9m��#�w���r�9\�������7q.���>A�1�flT��'��+/�s���ݟ6�Z�o�볓cm�.��#��OU"Ӕ�l��R���}q
b� �qNJ%6R@stt(����c��S	Jd���6���]�@X��;�� �J�cm�R5��Bˠ�5�S���Me��3F����(�*D~�ѻ�`�e)U"�k`�V�P�]9·G�Q�[�l�(٥�e-���ۃ
���({ף��n1�g�X��HM
�k�l3)�o�]�m�XL�Q�j�g�����\��E3K�u�2j�㶤���-���Y̫��zA5:v�����K��<�����_���c#�l�Z
��n�������{Ě� � '^�d�ȱ(��#�%���.����dT���C�l�����f(� ٠�kqAu�Bȹr�C��F���^��?L�ݒ!��;H�ut���x�3��!�7а�.���Q(VE&0oR��F:��cʰ�LN��H�X�9w1�_��%QjϘ�W��[9m�H��f��Z�Y��)��r�2��a��TK��44`�<M�s��f�A4v�xE��di�E��������y�x!:��`��ì�f�o���R˔;T{�'�_�-���T`�s�r9�Tn�!�0� 5�ߒ��_H� 龀�e�h������Q<�%�G�t��2znH���e"	����Z�<�/�����<��Z�`M�e_�OB^����/ޕ�k:%�m��^y���>Ȅ��DM���ÀM%�ұ��ʺ��>�[�'��cu�iAW�a���#.�������\�zy�!�U�e�u����;&�4��� �z�̧T���"_g�mA��魨m���)�tV������)Z/-���.���e�I��S����!� ���<g�7δ(S�H�k���@�����f�{豹�t\B8��!�������B:G�N��-6�-i��<��-� �J�0(Ǫ;�ڔ#q���g�&o�q���<t=��(�2m�뷺to�n�)�q뱡Μɦ�)��-T����jI�F��K�Ȉ�tܵ�]m/g#�] S'ߜs���'�5^�����F�K6 �tC��[��i�N�	�����)�=�_�f�	�00��L�_M#� ls�Hnt >�ݺ����	�.-I�|}#�d�|�U��*vQ��
!�qV��(�ľl����
.W-3~p,����E=�2�8����k�o �Mk&d1�ۥ������F\���
����F�J�tHѾ!��:�v4��3:� S� ��%���Y�ElM�y>������T�i�����J�l�/C�!�&���3�!V����&�[�� #=Z^jBC�Dp�RZ�� �嶢-c�ȁzܶ�k�nھW ��S<U�.��"�/r[5��Z���9�y�l�sc�� �.��ˇ��]к-��n;�Op����/lDF��Җ�y49�VB�c�eI�%kq��Sn)?��Ie����e
g�el����J��������nn�|ҳ���W��҅����5�(���0g���4("'Y�/�UP5��2#������'�T��ǪV��("���v"_z�C�豒 +$΂˘ru��1_H��*w*����O�I���>���*��l����PCs���(WyZ�܂=fMO��"3�M�S��Zs�;����c�v�Ag+���B���s�*T����r�~c�7ʑut��Ts�����𰛡�'�$*�Qy!�J�E콿�$�(���Z��]u�bQ<Ub��)ݦ�P
�[�ⵄP��9��� ������S�{�d9�VE��Rz�J��V���]�)���nH��7��`>�
�R��Z }L�{����a��;>	d<�V������<0���Ө����r�ك��?V7��H��[p��Wr
Bc�G�B���µ?G;���ăd�)B}��Q�ӹ�P��DH.���%щ*�#�[O�Ǳޫ�)��������澛]�����������*�:Tp��X����(A��i�~6mÊ7lB-�oH�v������$y�z��F��E P�[x)�KW�)��\C{�n��旁{�⚥�{�H05R��lgN�!l6��H�tAx7�F�h����>h)&�� �KM�j �5���QfN9���;=*��<������i�8�Piΰ�����Y��-$���Xu>|F>��Ty%�������Z$<d���Mw[��x���D�w2��[6�M�5�e��R�����~<����RB{�N��ҽ� zU]�1@z���z_x�p����u�\��@ྎʾɪV�e���bq�tuJL�$#¢���4���U�K>4�	��}�T�=υ�י��k��~A
u�n^I�$�B�qW�����k�#��h3����ɏ��TT%%��Z�2xV�S�ϟ���N\�O�j���$�%O��&������i�_ZCZ�I��}��)�[U��мj��l�Ny�o��PD��U������9c�DY:;aȼR�K�1+��J?A�ջ��v���?6�VB/��x��������� S��M�����<~|S"|YU��S��̀1"Ī1ʱpE���g]d�AO/�q�ai���
�!�n4`������]�ȥK�q��S?*S�$����i��r������RI��x���Z��x�(��� ��A�w����ǽ:��M��|%}������ېy:�{�<�{W_X�^��W%qO;��K��Nhgԫ�]�B�Mχ�Q#'^E�h{��m�L�?������\`59g6�C�H����_��q?߽��(�1dqm#�����Ҧ�>��ZK_k@�Fl��\:�nHl�޳^g��QRU"z�uzfyQt�[�*Ʉ�m��1a��ה����H�}�0*f�_9���nn��h��
ң4��ZՔ� X�X�_�mb��fYx�>���x�_7�;귲���,��������
Px�X�?�J�������MqP:?���"��j����ʫ�E�����($t؊��@!/fxI�2G�yG|U�
Z��Si��^;�p���s��2/U�]/��G�?Ȅ���v4Y9>�e~��e8�u6C��İl��K�ܿ��1޲u�z"1=3h�Ȓ8v��H'<��IA@ƥA��G�re�E.��s�F<%��R��:Ͳ*髄KC�g����2mem�񧝤�=��iY�����l�5��.t
�Dӌp�_A�V
��"zޘ�D�6�I�+e��n��ٗ�<���QF�|�Ԃ���{1�I ��I}��i��E12q�wh��1+����c�+����<�Yw�^Ы���H@M-:�O���|��kW�#}A��� @6�'�jU��d�S���-�ޱ�&҃��L9;�[��ܲ�'���UC+�R,˒��	�":u�Gc&-��zo۝�v�M��LY�'��·V���1)�T�"��x����!̓0K�&Q�?����|�ZOt4��?h9Ԫ����Рh]o�M�|+�_�^�Q#|�,�<��e,b��ɗ��-�lI��i��HP(�-�e���5Rdq�-��3�«#0��;�)V��K�K�J+�?\�˛$��a���h��2��w�����S5/�_� �|j�չy����ʶS:��#���^OH�"���ʣ��n�FG���n{�bE�/5ώSO�u~��R9�&4!~)��{Λ�(A,����s椟=�
�?��?w��tCt���8��41�?��(Z������־z|�Y�_�Q`i�r2������L/H'�g��
���5�xo�`�H�������X�X<���K��G x���}��/!��'��z�i��q1�VW�;iޞt�6�,�w��:X�yjI��]�~T̠�̩��a��!����e��^���o'���B��V�(bc�C�	��+�wTw�!�m����nF)�Sf��8e+��'D��G)���2Q .!�N���f��^����h�Ř�O3��YJ��_�j�T��l�O��YS���\P�y����Q�.�uG(l�z�Cz����W�?~E�`x:S���֭d5��\2�\��Ev��A��	C-��
�ˇt�%tzǀn�=h�a��W��h.��1�2���� �#s�+X�<��mm�0�B����I�>t�_mm� ��M����9����/�G��|�*k�㦌H���-�y�#��Q���dl�;��z��R�G4��>�0���f�2=��S|/��Cx���J��K6�L���Y���X��*X̍��p���&�M��K �]1���5��y�}�gXA8��N�bm�K������t���D������!ւd���XN�@,}���r�V��ɦף���p���J)$����*�u4o���.Vng�4gL��3��j�#S��+��5�!jv�#�t��V��8b�"�;��W2w�G�l��N=ه�f;\�ߍ%��	mW] �J!���r��Px5R�*�y���,����r��W�\u-�~��i! X\&�P��[Ee��	x,�Փ�{WI�/:����\��'W�
2�a��s
�~��]ߎ��϶���=*DpI쏤t��k���	g��-�t��}�r�o��E��߻7��)OTu�!��Jh�$�2�����1�j���`�^R޲%�k��ǅ4B� �@�=U3�&�QL��/����4��dbj�r}�������scSVKf��lJá�����Q��)������J�o^]�������H��*��8 t���yw�Pm8:px�r~:�=x(3|�|��⤎�h��X�Q�4�琤Eօ& �y�3��(�wC�ڑ�|�G/�\G�
"p��|�;%�b�Q��D���.�U�z#�U!o��6�B��h�$8��jm���2����݁��Ֆ��0!z�0W�t˼�|[�v;�V7�~�[�WP�E�O��Z:��ۿ�C@�'�O����J��*�\��q�~�6�� �����C��$�yۦ�_J���|6�S��/,7�iw����3��ȏp��,��]IS�O���q�b7�[�M����Q@l�o0��/�3T=����ƅ��vg��G�W������/�U�'Z�dSh�.�Q�m8<`�m�f�&�B�y�V���3��O�5`�0�F�p	�'��߇���::)r�����w�0�A�G�u.�z!d�VTJd�}�'��\d4e��qNt &���c�BO��	k��e��An����r!�):�Q�N����؃,���H]�O/�m,�dv�k���Z��r@QK���URX�8�>O4����ED~!4�Jl#��FnǼ�gm�	�ʰ9�4�&EF!{i7p��q�����{�ᅇ��o3�?ē���_<�p ���o�;F_<>�.�_?��r��.���?���B�B&-X�\(��z��Y�:Me��3NK��Q�!�$��z��'��k��N��^�%��?z&����B��#�E��M^�Y5����JO��_�9��Yy�(��UP��j���BL�-�1�A�~J?�I�Y{ՕA��i�dOA�G�BEUΛ�WE�T�{��P	�R��ٴ�>x��n��D�^�YC5*�#ASd���{�9�	ar�ڪ"S��j�ᡙg�0��\h����{^%��5f�p��lb94w�^kb��BȬ��dE�g���r |�t�NH�����&���-�v
rQ�x�0^��mK����U����)��26����7�T���Ɵl�3OM�LK�72�g��B�`h�aY�������T-���ѤUdl��wU?�I�iв�(`�~��� ���JBB���.��WÎ=ā����<3��=u��y>8����P�X}>(
=���3�}�2��=`�X��k_��[�3ӿe������P�Ţɻ��F� �H �&;�-FU�@��A>�慕{����Μlڐ�'Ü����O�G��ҒkE�����W0��0��Zӗ�2T��XH����O�[����.C��8k+?���u���0�ljnZ�I���v&�����b����3���!s��)!�X�1`U��+��o�(o:�>�y�[�Z�w�z�]^l�>�g��"�w|H	��}�31�.'8ۉ��䟢gS(�c¨��e�����l���D,�`�OLu�Bo�r�a���k3 �$2}}��L�dBx��]&�_��c���w�A����ὲv�nU����ҩ&���,c�7.'^k��
�����(zDQEhA
����6a�~�~j��D�^���Y�o�H�!}�d�g�10);n�Ĳ�Jq�	��;$���]^ϫ��2��߈|���Ρ�5_��b�Ώ�t�M-v<'S.z��q/�\�<1���ZY�6g�߬<
Z��{��y�*�Y��c1��C+U����|j�!�Hl$h��ۻ�ð3%[2Z�t,���a�-��'#ǁ׸�s̈�;���Q{u'�L�L�'ꚯ���b����
�T̌,� ��E��s�f\A�xV����`�B4\�\��C�B���B�*�n5��U\��eb����S�b3�|�y�X�.�I菏^��	v�V{p����ho��P�*�L]~|`g��fI,��ˇ�����H����^Wa�G�-��[�`J$W�_
����Tf�۷q.C)=
l�x'��x�AV݁�}���q\.n#ߒcGr?�]�U��ʶ��7�V�%�Ppb�<���HYh�w�^|&��v`�ȇE��I�gk/�M���"�K �-�Z��E����$s�W���Xr���HEq
�;�@��-�Ff{�ͥ��s,���]z�������Dt��Wqb�z��eI�(Z=B�B��<0���������a�7�� ߱S�p�CmK+.^�Pphs��\wR�ه�!G�R�Pn���+q{��0�F�5ԥ+&;��l��)s���_Z��a�ld��Yt��C�|��3�qR<.ih�v��x��!��4�c��2��mP��t��zc-f�4� �)q0^GR&*M�