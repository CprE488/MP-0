XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��7`����H���T�
����8fp�s&��36�A	,���|�P�0�F.eu����C������	t��8Q6�K���x��d>
 �qK�[YJ��Ԗx�;N3mVV�uGIM0��kk�V��_��_6�W��ǅݤ<�Z��4F��rJP{�'��uY��3i8��z�D�!)Q�������&3��7����~�;��s��� s�&Uo:�l)=�m��,y���'���;x�/	�^�M��L͞��;t���8Ű���Y�]6|�^EʲB�
5�n���aj��f���'�oPE$��w���w���w��8�T_x�.s�� �ͩ�	]>R8�$}�7�1���q��g�f���=v�8�;�Y��6^_C�~1<�����\o���$���\��z���!A��%�E��*�;/l�bj�'��ڒ�^���6C~���4��}(>٨ϞV�ߢ���6�-�
��ڟ�\j<W����8y�i�CMp�R�W6`H�G��*���Lx��"��>�oҙ�s ]p����A2X6	P�C��IC�� sT�,�M��O2Kx�F��Q��iS��`���)��}>r_������x�0U@�ϱ��;��%22]���`�V��~�J�� ��z��O�h/r�PZ|��%�Y\��d���҇S���?�2fFC�-e������^����|�
���J�d0@�;F�U���-�� �^�;��*�HӚ��]� �������T��-�~�?T�]GJ��t�XlxVHYEB    1853     810�s����=����+*�6��J�2I�-Mez�"ۜ�~l��!9t�]�&� ?5�ii�� �i���Oc莘�5��x��!���䯗ǲ孼֍�'�l𙍙��e$����j>�T7�C4p���y=%��Ĺ��K���$h�V��b�6��!ߗ ,^ob��\�a꒩�Agg�P�FJ)�iӸ8��ـ	�R�u�5�D�!�%�0��?�\�?��8V����W F�]�����,mLe�/�n���cE�q�@���)�+�������ߡ6v$c��<�Y�Sg�1E?[��E��K�Yt`3� �B&n��eC� �v(�����@�
Jѯ��.X /&Z�+{�1�%��vB��r���L�ؗ������� "qA�Q{����~i�����Z�`��� %�K���[`R�
x?l��k��{<<4�<u�X�����>�����ܝ	��9?�c�P�޵�R)�$ԃ�D��k�a���_�^y���X@Xͽr��q��̉ <eC;sN�����A�h��x���e*�`>NޤV甿uP��8��NyHE�wȤ���>�K����I��|����`��h���J��Lv��[%ya#|#��\�kC�|H{�V�Ɏ�ZT��[�G����E	[k��Ȩ@�dY��Uq��w!p���^l�z�?�F��ě\�L�����ĪOet�k���*�k2���{~��$ ��?�� �����t�C6'��Jw�6W�����'���
~��A�VK�cia�|��z[����y6YY�7��h�������+k:e�;W�a�_�u�Ϋ�\�}8�Z��F���v�peR
�� ?@^b�J �y���j�xl�)�d	�$G�q��\7�Y�X���Ԣ��ڥ��O��{τjhw���	�+�DH�٫�R����-���$*0=��5��g0'D����潃��6|��ʏ�}�i����Gkh�3G%}�� �!\#�NQS�㲚|'����؀�;�~�؉c>�>@�t�t�����C�����V^�m�6q�����d�ң�lRp��hU�:5��찤 �G<{�X���K��I�:�d6&el˒��JN�%p�Ģq@,�,��M?H҅�Β�\���P��+�/;��p�Rt�4H�Q�;�T�?�z9�kv+7Mh�@ΪW��K��w�^��'oOa�B�����a�#��qQ��� k���Hl��k[\�������]�>1���e�E��J����C#�������}�*YNd�Ҩ��
4�Qm}
r3I��χ)�ш�A��a٧Uk@I�t�)���{��J~���e;"YF���($N,Z#<����%pӵ�^���qC?o���
hu��cI�1r5��VIn��AI�����;�_ނ$�`���-[�2���)H�3l��+e`y�O>�b�I��V}ܪl!�%L��3j�1c�/JQ3��B������amє�5C�͡�Q�J�4��f0ba�u3��b�eS�Ct�_��W�K�h����Vx
m�J�v��X)48msH'�Q}c���"5�A���Z��$
R��V��"YU������JRp�d�C�4�NOtD�y6G�\�Y "�O��﬈�W��T�J�Ei�w��NQ�_kOg�.����	+7�{v#�ۣ0��h��O�=�3�'��`�`|W+�FeK��*~�(��a��?��4��%�5s�!}�Ð�yf:Z�篾�9[�u���I[�?���k�]բ�E&��Zsk��6�q�h�%��<�#�Ȧ=D�:a
B�A��:t7P<<-$=!�T�:Y B�8�I�M���j��F �2.������=�=�L��4�q�u�@������^����5�hՓR���\�W�%tz�HV������Zxۗ�:�N��L݄�����.�J�G���p0���-��H�{�u&��3i�;�/�S���a���Sr��!`l"ؿK'��nZ��a
 9H(?w�8Q�	(���(�1�2�s4U��6Ivd�!i�b�8����<˂���I¸�����Hҽn��A�CKNm/Rҡ