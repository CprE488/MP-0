XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ZH�8��y�m<^ޣ�Z^��uU����]�e����(]���*A�"^�>�(�g�ЍI��f �2��CD6��o���M�S#7��Y�.דA6e�@�$��۶]&���z�Fc��森m��u>4�H��%��4K����\��}���J�a��X�]�*w�R�����@��@�ƫ� �"Q��w��>a|W!�9~E�%S�҉% 	�L ��i�w5,�� �b�Lݛ���둯dY*���Y0筑}uJ�M�?�?��4
M�9��N�cY���%!a,�i"�\,�Q��გ�-�ܘ ؇���~p}n�B�B�"�΃�75X�����'쭱��_���"�����4��r p��5���ޞ��p����S���KҒ}�~X3���FV�0�^���5��O���¶,������������1�_]6ݳ%g$�(^? v��A�y��S����9�X���.�\��>���x���əx��퉐Q�:~��M��̗d�{��U����h���̮�#��'��sև�3��w�w*>�F���R�U���7�RNw��ԏn����n��W�ݘ
Z���+�2�K*���UNAJa��=s'v�o�@D�s[�u����&�=�=��+����z
 J�b�at�kc�~��K}�ߗ;,V��/Oii�\���� \�iA�b�j�'��b�Xh�4V7b�m�+��9��}�C�돃�=U�̀<H)1��h1v q|�\XlxVHYEB    dd8f    2160f�u���Y�u�^ㄊǒf"�C6���<~{���q[��3���4�7��j� 9kd��j�� o�`����mVZH$�R<;PL�|�"ăJ�+ؑ�WR�P˾�dݮ� s���¦d�e���AP]f$lE�~S�:2M,�#��vNK��oF��r���
�j�+z@,c0U�*B�����8a��C;�W�Ƥ-} $VGŋC�m)�	2�OQ>��鍇�8i4��>jL�0iZ��^~\�U�p���" ��P@�ҙk�#��{*�. B�'�E��7�s�����%��f��>����:+q�P�V�Ф�}�������ޣ����:
#I�����+4�r�W*߁o4rARG�+@3h�ݵ��R'f��x��C��A̻}�(��
�]���?S�[d�)����d�Rp�W��)��Tv��m�=%q.Z���(۷N�2yT^:f���0Z�"B��D��d=�4��ׄ�B�ϒp+3�ּ����RQ��ρ��ʻب��Cσ3)Q�����3�X�I&�q�}c+Te��oH%�����z�� �/�jD���n�}�p�@�a1j�t.��P��S��5����k���C%���z�
g���,�����0���.���b�xvgЎ=#d��Փ��~	J���T���'�z������RL��R���A��d0�&� ��@�`x�B�&�Jim$ʙ�5��������MwG��c=�����I�LC��bbB'$HjAr���ѽ�Bf?~�j�y���lׅ��@�_�T*0�N���a�w.Rއ�� ,+�5����:zˤ���h��I�]INsĴ�G��l��[�鉜�/�X8�Z8�rLc����Rv�o�_�|��jP3�֍�C$-Pq�B$�ts���-�]jcG��#�W��ǭ���SPZ��jr��c9�/�v�ꂄ��a�/p�/����������D{<�M@6�\��K�#+T��:6<�60���Org��0>�G��D?�n�VR)�=8	X観�U�݄���3��"�����W�^��2��LC���GΡ�T��g{b�w*|�:X6�l-Dq�7����I%��#�s��@_L��\�I�{9��7���p�l�f��)���zL�l�v^/vd����=�����T���xo��̭�}�n�Rk8������{��zjB�xJ�{�6�r-�T;���V�]8'C�?2�񃾁��7�A{��WŃ�|�ѧJD0F��!�C�0��	{�&�` �#|Db���!��}�Nk������;w=l�C�5G�ԩ2��j�� 3QH���PǰFnB�aI�i�u�p�b�2Re�:�T�~S�(�1)��&�1��m��r.%��^�mq���6�{�u:��()$f��ٻ��ފ�����$������ZQ�|M�W�ɧEle�Wce�,��Ι�Vj);A�	��[9��lq�� <�{�BZ��d�����L�T��Ƒȇj
�G�g���GYj�X����j�d�旼��z����tPG�_�^x0�>�����b�AU9��p�"���y_+�ːc���r ���`.;�`�ԝ_��|�%�p����g���N�^�	��=��������t�H=�n>�A��>�oơt;�;z��3d�冤�="� f��Ir��z_:�Ȕb�aRF�]jc5 *Ru����{$��k�8��˳ �84Cg)Ư�$�Ӷi野�y�o��f�������$Jf�6��Z��&�A�!و�o|�W�9{ԝ����r��b
��h�ܼ�R���:�
P�͡����T�M#*I�[Q����(u����j�0���Ȗ���'E������B��!��50��������/ �9.�{�!�>\�\�C��䨟���;~PTei�d�®O��3����[u��V��Q,�bn�~�˺]I�"w�(
^��G�@���S2�M���KCĪ�lT��/�4?2V�^Wk��8s���}�	ȩQ��
����}J!���Hv	2~"3Xe����y��޳'�L�_+���k9����Y� G����/ss�3/dHׄ��e.!��w��.1�z<J��B�@@t)��B ,,�!���ǀ'�ז��R5��b�������g��ŏ�c������c��:�Y�!$�������F���q-���C���
��h�݅a&��}�S��_�XA��I�0ÍU%��*�*/*O7O�Y���	Z�1��]�+����߯Q��(�T.�� ��_��{G����V�%��oCm���3��m��\9�&��>{�2���V�tb� �RSEߝш/�`��e��p�tJ�C!hvV�*9�^0rd��C�#3�n��%�8R0޼�꿃�3M��MlQI�~�8M$��{%��~ġ4����l���ԍ�8����p�
�~��~�d�j��'ɀĽg@w�&�U�~�&�������Y�P8�~X�d�������vm�|�rk�R�j݋�x�C�SE$�@N19L�Q��ûP>�Z�4��.��
��<bk>��.9;q,���&m��!/�lº�?U�Įh������'��vѝ1�]�7�[b�N58[W	�6=6�Id��̰�u�Ԕ����{��>jq��c�H�!,P���>1T��ă`�N3�@����h����t���E��q.`j�?���"�L%����#��]�vw��a?&{�=Sn�L��q�E�B��:W2�Y�����յC�:w��ե���ӽ�-���L˗$"@M�.+,�]7C<a2�q'��c�ݖJ�U�<U����F������U�`�呂?GF��޹e��:��;��2��2�,��K�e���%�m��q��P�8[R
l+2�4���Gc�u�q2��ބ��]��C5ۯ�6?6x@\��	�yש�$ӛ��֍$Ld����4�Ti'?��R�D-�1��q�`~��pc��@&�_�����m�x�5|���K�)�j^{�m\�Mďd��B���;X�`S���_̈́KѼ4�x��j�pn�6�a�D��1�6��A��6�5�����z� y)��H{_��.�[He�_f*�j`�S�[eZҡ U�8g�74]�J[��\��%��ʴ�H�gg�����I'�<~MeI��R�?"�k�ˣ��D�C;�3�R�s��v��	���Z�ݧ||U*bz[;�DW���m,���S껹)d��A�prV�,Ȇ�"Tq��s�����Ax��G��f��ptf�Az{]���vT��i+p֒K��B@��4���`&��"$�[����+�1�A�)��ʷ�6�<�ǲt�[�J�DXH&�Dn�/Y�V��RM����=�꡻ȣ[w�K�vNƆ�(���Q%],I���rO���Z� $�3�����^U��j	�4|������v�}���ďP
#��!�jj"%nLM���o#���/P���=��H1�%2�|�������A�9���F�P{�������F��^�{�שg�t����B1�%�e��MTw�5䮺��b.�'�f��%�l9Ws�3��%�^�5�zSa�p�t6]�*�B1觞)�;�sP_Ԗ�����}�� N{C��&8)�k�j���T�@g�d�9�s��)m�ʷ3r�3�=�;@�{��q�z�����ztŔNH��"6��s)S|�b�C��x�v,>���J���-ƪ9cnSX��D����	�D\_�(A(��
�잊b���ß�D��D�|GŊ��^U¬7��Ƽ��%	�d���10��P�
��I��a��Tw�I��\kҌC�����Lo�
�I؂�o�#�!L�;����yOo]��/�QT*Ӌ�M;'?�*>���o�V�ʣ�_�֫�g�����S��Ǚa�zB�!����V�`!�����z�8b��!Z���xN�����)ʧ��p��3���3j��	�C�?�P(9L�7���;E�"�0�qDD'+�x�Z"Z�u��<h�Z�b���F` ���툮�q%��� v�ɔ}�� ��!C��P�a���͏ś�t��!)�zfk��_�&�t�����W0RLô���M9�A���1��$�R>�k���lg�yy|�
:
��B���GW�N�bt{D�ȭ2s�؝��w�&a`�s�؜o6G�@7r�'�&=����;�,.��$ �9^�&��L>�E(@�ax~~\6�[�:���AYd+���,�K�P?5��gB+}=���D�'h���<'ـL�ם[@��e�������a4k��>��m3��^W�("�`�!ڮ�[C�(���W^�-�!�N#�k�H�f���!C�HLY��=���� G�KlB�WV���z�c�H�3�ǵM	9!1�$��v����`�$����.�ag�`nl0�ˢ���w����鼭[e�� �gC���Τ���q`fQ�n;DJ]p_Ã�Lx+s>���� N�_U	T���������+��d���fM{��}�UD��x�U��%��O���j����e@�&?�[��.5�Qל�}Lז
2l�Q/󧜁3\�����NÖ����M���c�����4û��`�Z~�e44.�B �yW�s��m�R����	s!��O�|'ሔ��i����{+|��/l&�n��Z�1���k�Y��хgk7��[ya�POEWp+����m�#����}�~�������N�$Y�nۡ���~�A�c�A��R8���g�ܸG�4�z��3aQ����;�\�%��Oϑ��aS�~�qb݅vb�QH;7�>�̉���F���t#�/�G�u��͋�Lg�%-%�E� ��J$a����2w�[Wq0Z�q��cn�"�T�k琺|��>|.�ϗ<7F�)�y�c�~�
�l^=S�Ę�v-��c��U=�6f���[��X0V��-B�����Y��&�Xˁg0V���#Ä&{�kc�*Lpa/]�)e�P^��(�V��D����X�����v�{� 1P#PX��b]iT
�\j��Q�Bѽ:N��^� n��(�����q8�Xi!���g�j���i~V�8���(�W7�6b�r5#���-���2_ӽ��|�-�Z��m�"��Z(H�!�����6��En�S�v�N���>߽�c�ǝQ���Z,�?������˞�̦ʞ�W/��&�J,TFҭ*gȵ*3~�8`���?i����N<�(����LƝQ=��*!��sU��y���(��10�3L@�-i+QW.�4�*�;S��~�H�XV�&�b�Z�=Ou�I	���Dcȋ�Į�_�n��- �l��	�����دi��Z��\�C�+덱˯Ye��!T��麱.�O�������z�z�C&��z�3O�>�P7HF[ȿ�Ejte��Q�$�Ćj�g��	?�Yz~�.�fG�Ǒ?O�F�.Y���1�:(�;c��9�y^�&���bN&�w7c7xt��q5d���n��Hs���BƝcn�[Ӓ�m6<�.����b6�#�϶�:5+�����g�������/�ڍ�e���r�i�|�0&����U���=�w7퀡$�"KoZ�5늗�ݼc�7�+[\>5.�r�6��'�sr��ؼUwk��Ld�h��,%�,�:����\!Ϧ�c�	iI!7��̅N)��ܙcp��0[��6A�l��Hߓ��g#׵ ��+`�gY�k/����/��κ����bB��D���IW�O�D���Ot��t�n�5f��z�+�g���H{~�S:�[���q��z�sq��7��=�]fp��H5Y_Tv�����%��ͷŮI/%ߥ�nx�H�Eq��4�8��:�SǔV�.W�ߤ���V���{��p�����K~N�!b��gr_vÞ�֠�ܮ�$�ٺ��q��|s�?���Bʮ���L1VHu���)�9��<$������"fV[�2�e؁̷I�ZJ�ؚ^��l~{�~
�������o��c��fn��lvg����3�M�n��r4��W]�G��"]ǃ��u�?�E�QJ~�IQ�N~�(
Dے�г�t6�W=�tF�f#Lwp����j�Ɩ�Jp�i��P�%E�A��J����1�+��s��Ѣ����x(�Z���
��&5�o��^cp��j~���]#���`���g|j�#���X㈆���i�=/kǓw�Ii���nU����&E��5"�mV��F�Vw�(�4ę��I9�ef�J:ӌ��*Ů?B4��G�N@֫�D ���[�q@��~�l)^ظi,s^�3-+w8B�dI���G�C�(N�5׊2*m��2I�<'BUθ��V(��S5ä�ǟI�&��F���ń��p��������bV� P���q���B��/Pϙ���)�ð�$z�6��E��F�@�$ٝ-�),9vE�h����ɟ�N�Xr1�*R�"9%������� '%��tE*�&�8���ɟ��L}���n�{C&��_=�����.E��1��+�yE%��{�Hu�!��/
@X�eX�Kȶ�[ۓ���+.�ȯe'm=}�����jv�
�J�P��;z����{id�����ǎ,~���fFLZ��,u�[�$�}�s;��ο�X�w���y$�Uq�UІ㏂:I�/_e�V�&����E��I8sbDe6� �c{���
���d�_%�}���q�U[�{O��l�����k�	z ;��7�+]��V����u-��E��b��.b ���;�t|�'cQ><"��+����0;1�?3^�&�m#ddY��2|����ݺGQ��(4����l2���<M�>9б�y��.�@�R O�,4�������4�6�B�g���\5��C������p���_T%�s�^Rʹ���I;b9R���O����TQ�.�[+��w�A�ͱ�l����R���a���;��p�k�ɍ԰�n��CE�D�Dj��#aC`n�ܘ�Ib�'�-����]H��Ѷ��l|bd�Ӌ����4�9Y,ؿ�6EC��ԏ�%����`�|�Ux�ĳ��5	 m�ϧEǆ��ϼ���#հ�~a��h��վ4��,�v(Jp:�ѽ`G�X<�.ML�>Sƿ�H���8�N'7����"H�-XE/�*y�;)�o��M�����y���P����k�Z[���4i7'ڠƑF#l�/OI�l �!��7{��$�ȝ4��c|Z�'�*�V^E��#1�:/��-���H�We��HH�0ɟ���^�Ж+�T�����B��(Gܹ^��)��.22w<�ψ�_��b��H���\{������^�g�5�9¡� �� Kfovu0�q!i�%��0v���z�TV@��X�^�+C`�@_����Ax�8��@���g�� ?[+��h���2��X3Z��NY�m���͔�j�m�[y�Y\��I'd��9J�ImŴ�����ĝ�^��_��'d���p,��2�0�I�x-{q~(�!�{vy��܎��Td���9�N�|6j���"ծ)������ݦ��z�'���*h2L���.-ZA��~k��?�C4 �.��^�>�3��t��x�Y����3��X߷��k@#�>
��8��5��ʧB&+��4���dY�������ԩ����@fQ"-���g�q��R��iX��Y/]�=K��͗�cutH%�_���:I˂%3�l\���HqyFu��)p-�=MS(��F'�FE���� 6���,�p9z�z7K[��PT�a�����Y�8��;�X3	YWW)Xm  a�֤�{���!B�BsU��.\���Kt �H[���h���I<��j�V��?�o�h
���W��ÛF1 �S9��Ӏ��r
#�i��y*�ͤr��/����o,b(Fd/r� ���C��4��;��$^+���5K�V1��g$N��Q�/�����^���`e�����-�h>���a���s��,�T���_���:X?&����bо����֌��f���&u(�l��x�Ӭ�V騦�x7�fz�a����o�5������5��طNVMƤ�{2/
�iM}��~j~����o�p��A�T�5?YP ��p���@1�5*�� C�H;P=k0P��y�v!9�%��9���^4X�"u~B��;5�^��?t,�����^F���~��}��r�yMJ5�E[Y����a����$W�N��ʜ�4�볝q}�Gԍ�7`k���%Q�4P�!��%LD<0�ew���Ĵ>���n�w%��S�_4G�z�r�%ZxX��t%�������$���8��jX�!믧eG��5�UI�@�.�uЋ�@j��=FH%d���`��lN��.5�B�,��r��ɶL�I���.��>nΑ�EtBC�����.