XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��hKn�_v�ۉ�Iz������KI�����kW�Γ�L���?�^tĪ˃m'�m��E+�$]'b���X�"�������TIge�Õ�W9����Z�o6�&o�.��X����^b'
I��Z3ؚx<7_�3ZnG�W�R{�~���b�uGo�B'�Q�v#�8-%x݇�Emx�+�����t�_B�I��AK�Rx��Ak�1���%�lWو�7xؘ�ï�n�qR ��CN��lp��T8�we��Kď��Ƥ)�ki�*2�EV����,Pq�M�|\�@�K���UӒq.��N�M%a-�ͤ[�c�:N���Åc��e3��2!&�n9�ȰƮ�$���`s9�%�H�wd�}z{��LkiWQx��ue�6ހ�'�V̖C`NAH�-��rdB~*�2�����Ԃ���%sҖFe��h�I�f�R���O,���nN�Ru-�� �xd�~�\��loj��&�#�q��FC�rL�����Mӝꑼ���J��Tk����WB88�qh̹e�:��.������r{{���B%��=;�y���Q2m'n�dL�10 ��9�'ϵ���S.&�J��G���yX�p�k��h��?�^t7�`������FND�=s'}�ŲHZ��DGd�o'�oD��w�Uj��R��-��N�Ρl/c4�?>�C�Ep�O���]��'��[�]s+��s��1d��u�٠���3�AY�|ؖ��Ob	� �.|j�2	F��c�a��ې�.K�	�XlxVHYEB    fa00    2040U�c��6)�0N�����9�{o�|�c39(�G,������s� 9
���!do�\���ڑ|���βw�v}���V��E�/o� �80 )�8Vhڊo=��F����(�Y�?��hm��b���.SR��V?	*��i!����5(+=�B��e��Y���B~��KΌ����)�+���x$[,��C���u"�z���&���ݒ=�*P���ݻ�"j�KS�
�^��,�U���\п� �ǄT�^��b�79�����Z0C���� |�^��Ese��@����;�9��保,��Kg.jۮ7�Σ��|������d(�etc��}��pɰ�Ӹ�ۻ<��S�\b�o�T�M�7��
�~�6p��;aOP�^�1����WR���!��ȗ%Z�zC���Cz���i�SU 8�Z8�1Ög��+Q>đ�{3$]�����^L�X9��p`�d6�.�+����y	�B?k�ꘓީQH�|��U��΃��i���	�L~�M�ˇ*c�ۇ$I�z�H��d/�a�ſ��}<��=�5�<DƊ���� x�W�X`�g�q��Z�Vќkk�FC���:����bPf��yϜ��E�D4��{�J��ά���aF����arX��Up�Ԍ�(M3S;SVӀ��Ý�3���0��`��~�D�=�4���+���kW�g]}}���g��Y+�?�ВtrY�ރfi ��Ү�p0&V�q���b&Cv�D]$�i�Y�Q��ay��X̉e�%5B�R�T�����N?�?@��#�n^H"�9��9�U����aJ�y5!B=�|�dn���E�i��v�.������(qZl�D$�"�Bۃ�3��oB��qt̯��v��y7pH.]��~�V]L\5��Gܽ��M�ʣ��?��d��@[��?)�xX�դ݁����`�ɣ�`6�D:��7H����j�����K�J�X(ttǹ[�:�-;M�b��xi�-�.\�:x��r8c�a�s��|w4��qem|`�LÙR?��w��ϣ�OoR��-�����8��v8�:����x�]\�TX&��H�ޗ��4��{;}�����.�nk��?C��u/�e�s��x0��lC�(P����2 s���1�ܣ\�M��ö����y�B����^=�o����c!jW������"���qr�#�&E�)`+>&	�#%sB�R�_$�sڕ��'���N�]03�o�¹p��բ����ܑ�[ B�5������7�]hj�S�1&s�T}�f��m2ח��Q]ȓ�Z�6�a��9�4	x�����ε�g�@��(۰]�dY_���>z�[���˖�\�r����7>#��ewǿ������3�v%�y�X�{�̱mkI�`u����|Д�x��Nϝ/+p���Hokrp��`PX�����M�Y@��/�g���u�<���S�ֿ砸�K�Ɣi;<���]>�������
Z}�o\x̐\kp���RI���t�8���exC`Pٜ����v�A�F�|�B�#�$w�+�����;�ދ��!$F-K��Y���B�}{��՞&?Q�W��8��w�M���7��� �3mV]\�`���K���Ӵ4�#ve�4ɋw�\�zjDlъ�R�!%�S�ߖ��{����NDQa=�
�;�9���0K��6=�|��퓴�t�)^~� )�M�;e�?P�p?D}�"�J͓�[$��U�W�vi��)�6(Y�ͲI��0�)��@�\�M����Ǭ�h������,J#��k�!�p^��y�$E#�%QM�=� 8�}�1m�[2��.��q���%��ܢ��������}�P��6��+��i�w�c�L��ʤ�e����:,g�ɰ_�Α�c��GN�f�sn���6����e#~_߇kUcXa�rn/���~���p+��;7�t
Y�v.��qӼ����ƴe�Y��e�߄PX��j��gQm���5�׹��QG���;���T9��ćv���z��cssm�	��fr�tSH� ���T�I��>�=�x���>$�$��<`�ј��aɼ��5�+{��E���Hɡ�5��5�K��!�l4=�,];��8���5�/]�8U�Ym��D_4kf�ܣj
(NV<d���y�nN^��8��<0�f�.��:��$�B��Tr&�0���9�	��2M�K�w,%�sC��-���6(��L�H�W9�GX�F>�)p^�&�:�'�t񂾳o��缦(8uWFMYg;r��Ջ��*�f�$X'�@�K���SGr��:j_~��2�� c�W5\CN�YL��f9|��:1��)�+����b9�z���������SN�F��8�;��;�$/��hʭ~�Q ���'M��iZ�����/����cl��y~`��J�^I%*��&��߲u����:��M����~�,B^�L���_���T�(����`�T���E��j��;�cV1)�y4����|M��Ur��X =v���{�o���c�I95}|X��)���t�FwΪ�����<�$�qV0Q8u�U���C���Y3O��t����/�����
�6�YWP�� k�l����3���cL������Ηl|�r�Pg:�#�^� �����  %��B/������_�l��Ɲ�/�w�ED��)�.��%����)��!Ͼi�ݨ������2�@Ԕ�<�"��hʾt��s?�3R*�&.����~""KG�r��bu�T�W���Es�6��H��'����6���d�t_O.�ch`�O�K�����T�饛+��#6��EZ�/H7w;�;������IhRi}L��\"�!�h=�l8��Z�]j
�5W�f���:dN�����0q�����ϒk��H���*�e�r�@%�R��� ��Z_]�3h�W+'l{q���͔N��rNe��[|l�AJ@�S����t��3�yBǰ�_��0��]�.g�=��E�o�bD�F���kTy��7J1S1=�;\����� /a��A����t�$�o��t�!�W�()������p���^W1�nZ�9:b�����1��
����)��kC�">��Qj��1d��g�)A_b���_� _��۔�<TcL��@��9�:�9�\#u�P��Ȧ��`A��iB��?���ٹ*/�;�(�4���Cv���V�j�\<��2O���ak����ij(,6'���rm��a��n�X������j��#���+j"�(�o](�,�VY����<:���6ҷ�U$Z�H�j�"{����"1�\��!�����w@O�Rw1��ЁP����X��f[7��(�b�u+��R��mnN�-ĘG���N����X���m�g$�_�nUS�.i%.y�C�T�Ї�IXgS����dgo�tE,L+�Ŭ�z��#�� g튵�,�QM�c�,,�l9.�D�ak��C��J�ߺ=g���|��ܜ�rY�,�!�W[o�4����=t?��^6�B��`7=�ڲ'I�O�~O�!5�\�=8�q��c�n��2ed�K��-�l�o���."�w@Cwټⴄ�f�X�� ����1B�g�Ƙ��?�w1����K�9$��J��&��v�[	O�;��.>?aqLۣ[P��#�&�æ>��#V;y{���[��?����T�F���{l�����9!�X��I=�A'���2���Y�u)�؀�ށE�a��8g����
׫vG���U>m_wHRvTh��+DQ���`��<���k:1�u&��]��"K�Nx����]ȷ��X�9�������+]�6�G$(S'|�1)�q�
�����j�#���FL�I�g�c����J�}���T�N?�XE�ӨrHX
�z���i����{�x5�N��<��	V�
O�����N�� �
�S���eR�Sm����]<]*jl��6����D�U�+u#h��M��xr��9�����x�(���Cx�Ȗ�GX�S��2~����Q�#ԝ���7�Ky _���X8�m����@ם� %�c����Е��"*����ӷ�������;�at+q]��]�R�Z�n��O����Q#�r�q��?�F�:`׼�쁐���Y��|NT��6<8��"�
�FI��S7�s��6R	��.6���Y�W;�z�T+zs�kD���S8b�Gå}�����ʤ��c�Tg�[�s®-+�8����>��4�����o$�j��yиDa�NƦfq
v��ފ�*'�rQ������ ���mT���Wq�&|��L����[s�{4�t钸����s��?f���`�9��DӬ������@M��	>��qQ�w�:�X�d*��0����\l,F�mG��Q���&[���p�D��%]
V��E�fh�2�O5.i���b���m�4oL���
���p"9�Q��-u����t�.��o
[��2�;�����ZG����E݃2ݦ���0�[��`�;��f�β
����pn8��r�yn����Zi�N5G��������j*`o�^v񓊳�t�(fޟB7����<��}Z|��6�&L�$1����C9eZ.�,aua�val��3p���]t���J�L����-ZE��C�ƀm�����069�q����]V��+=��Ŭ��4w'���br����}�b9�?A9E���h� �r<�!�`2���	�f��v+/���s|Wp��j�Π{-f'��w�{�Y� ��h�����,��ER��lKp���rQ��CB(������v	ܦ��לɟ0��aQ�E��*�x\�B5��go���JxX`�ܾe�k��#�g��}�a��7��'�M��ɴ�Z��1�y�bW9(�n�s��M0�MA�4��80�ڧsF���$��QX/���cHw�@N+�Q�gw��-X=J6׸��.�s�Q�����A��x�f�ڬ|���,yc��i������?^��A>�(I�)
j:/�Eo��Y�e�+­O��':A��MJ��&nM�Lj*�?�G�[���R�<���{�7���[o�L��l��/3����V���"�<~��6�Z/��������m��`;���
^s��s�3��h��߫�H����N�R�����vNI���h�����l�ڏ�L:�yS����=����5���<	ۨX<�.�o/����һ��#���X�#8�|$���pe��l/���m�eǶ��Q�U��;��I����u��?jE	Գ�]�L�q(ox��}#���D:�ٟlͤ� w��B<��>Sp��wʛ%�Y1�>�b�b5��d�شj�D�V�ql".�BY�a`ly쪬�D���oJ6���z�k�^`�;Kh[��J`�gʕD;o�_JJO�p<�-sc�;�6�X�J1ƻ��o;мa7���Ɠ.�oa�o-����*�X0���R���ߒ���A�ؤ�+��z8
5}5p��K�������U#9�H���vja�c)�T�d[�����(��n9w�c�\����L���]��;LL`�	��O\6������΍��EFu���H }�J�H�J�ňi�Z9��_�0KFFU5�]"e�,���!�( p`��*c%h��aϸ7���Y`��-�Wq�dX�`0%���Zț�}��}X��4�^��w�-��}�h�)��� 8J�aX߻^�E�"�K��R����r,�����2<�����Cg�r��6�Zþ��n�y�-�
�s��/?ó�c´���f\�z�k5cc�V�L��wT�&��E[��h]�k)��Rd�Ò��fȘ�1\�^�nU=\���PAQ�t�w5��
b4D�:��	<#�Jwy(a���Ra�%������b�\���瀶od	k�W��/�}���� ����=l�����v�T^��A��'��;��e��
�#��[Vu��C���6�������#��%�=Y_�.Ub��S�o�T��vGE҄ޅQ��&p.�l62F3�k%)�RD���v4ق��jlN_&�˟h~�����ػ.AU��iZ8����v��`�zhl��j�e0�-�m�R}��香��լ�0�iKڢ��f=�5�ޗ'�Qj�30��ݶ~b��˂jTͰl��B�yu���L1Ԕ��B=���]u�dfC���\鳠?��j>0��e'{Y֒�/BwY����L�W;Xl�����j�������U%iq�d:U�F<3�IhM������7y�x= 59)�ϋ��D�R�T�!1ߩ[�#�*�+��հԱME�l[� �,91?�oZ�t�� y�M5���lwsk3OȒ�S,:SWk�ewD�e��C��oVy��I����
��
�"��=�1Ǉ}e����
���u�;__�{�7{gI�~0�m��ſ�+�<x�I�;�i�4Yf�\N]��~E�hߤ>M32�M��nkk�1��M��î]�
M�m�x��(���S���P����k\W�3*zU��QY_N�z��b��\��n�q%�pJXI+��n��v�I�c����}H��%�8@�`(�~[?��т3��\�Vk_�}�;�{T&ӛ�GL�H�Ê̒|��]z�Q6��MM���[������ .J}Y�,�2o)5���uA�v�5�ԏ�$����4�M�u����4	ݱ�N����1�b81J-��kn,W� �v&A�����)�͉R����,�# �%n!��,Q��ΗхW6U@�Q���R8.qb0�0�kFT�D��-�t�-����q�܏⬄���B�oxH��y�3�Yz�L�������-�We��v��q6�1�^�$�aT��?�gZ��y�`.Z�RE{��?TX����h\�����m_Ҫ7����q7����B>>�0��@:�F�y�ǟ!�L�:'|�S����A2&�:�v\]��X�muaDݫ�-/)�c����QӤa���1�G6
�/���AT�p�u��Nͅ���_S��Q��ۤ��a=U� 5��R��BB��)������KU��Y�8�r��V%1�qZ�wS��������#��Y�J�G�[����IHM�����	@� ��xp��ceR�i�"�*]���gSK_����1<�@�'o�(�r+�S����*��5<���ɱ	������P����j`Q����L�U���Y�,\)��v6d�u���9��4��G�X���<���<� .vO�$�T�����"P*YE0K�Y}!�G~/��"E~��S.��l^�.Z�����g�.�������e��2�j�a{(�K��a}!2���'M�v5Ot4E�P�zS�P�A�r��_c�-֛��f���z8����6��:��5��_:�/�*����X��]��_��/d�㳶��/��(��䮻���q /�r��IhJ��Ԑ��8��erAA/�17&�*QlZH��i��i�f]a�G�%e-Y�u��B!���":��HX�oj��1�k��t�/���T_�&
��J���Q��J&ad�"�G���r����X�+�iY��v�v��D�n���5�A��p �o*'j �����H��m�8�~��W�}���#��#�{�A���K]�ޗN��%E,L���婢"时�M3�{���<�uhN�2���c(�-���JӄD$Ɩ�[�-��a2*u��@uR�EW&ݸA8HYlm��FB�LFQ3��D� �h���!���IO�B����'�838#���>���ku�A�i��)8_۶~�1�=��$�� ?H���݀�]��}�{�s�(gmb�iV �'�9��(`�@/����p�VU��.��_�3�3d�wm
�������jM3e��<�ĊV^�
����R^�)-��I���2�>��[�Z�,������̔K���1;����U5��B��Ǳ��fDz�w �z3 l��;ݪvץ0p�0�Vd��2ϑǎo�	|��	�y��$dnt}MI?��m��lt13��=�����^$-�ʖ=9�"�)g�q���jQ��}�$�R�y�6����`"ܐ9	���A�`kB�a_]��Hx!��]�pܐN�s(+@��=���0�G0�Xb�/\EVk<�*��+"Eq�;�mt�7�ӑ-,4�]4U|�P$��R�ߠM��qXlxVHYEB    4f62     b509�CI���p�g���Q7߅`��O��hzZGF���[��T�1#SܔSE���$�D��G���̨?u�Q�.#���_L���G�G;S�;E�X�8y��6�<9�6#��~�� TA=��ۘ%(ǘ�tc2b7V��KKH��s�e���B\\��$���5���u��n�V�!�8�=���'�1���!��i>rh�w4>~���=�&��b"�a!{�hF��V��vߣ�@�ʃ~�������{�Ȱ+��f�CH²,���2h�!�Y�<� c��`@ק�T�_`��(�dw����W� ߗY��J�D.�/"�դ���V��?�
����.0ʦ��텄���4��:�S����nebɆ�P�L������ڥS�Y�1�p�7/l!&J_i�2؎�[�x�A�����:��1�֥�[ȶ��n ɘ���nF�eYeqzȷRW�P�%��.�A7u��O+�@��_D�aca�9,��THLɧ�e{��來�H����%�����A��`��p93-�N�U��og�������6����	p�i	�R�fx����P_�G̨`�o�0���?�U�9hk��ɸS�&*�pˌ�h+���d�t#y甾��YX��1�|�ǃBSh,)9E�u�(�B���=�A�,k��C����qã���V�&��v5w��f�5�SƘC�B���J{)
�X�������Cy���z��	�=)
M
#��7��F�O�C�3��
���M�/׋YаKT�S�hHV��tS�E���v�aA����> o�&�Ȅ�&P����&Е{Y��BȀ.��8��cEɈN#��Vٗ�����6�%�C�F��<�*7�YJ�t��V��+�%��k�ڤ�<ϡW�Qn&��}u[fS�b�����(5�6@#T��	3�TǦ
�ap*<��;}�Y�x����L�	��ɭ��r��i���Z��;�xγ�����ΤgS��*Y��$B������uy�ECxZ,B��b�s���L�m'��9#Ý{�4~O���H̹�>����)޲r����4��;��n�NѧLG�odH�lh �P�oI9?��IR*4�J?�����DN�r2<�눽�M��Z؆kG��{�O�l
��_,�RE%O"np��Ǯ츪� -�j�@�;8���l��&� r����7�>�NY22y@+`l����_�~A`#�\���e���Ӳi��"����5�	������s��G=Zr��:��q$��T���x)jNL!|�Vc�u��%+��)���q�:���/b_jf�q^�ɟ�c��G�!9� a@�����PTRKv��h��pn��$�|��K��t>�Y�8g��S��L,���7�#�tt����U��`�g �S~���ڌ�R�<%�5c��{V�0�}	�#a�mi��3�{�J*�]J7nM���f��j%	У8A�GM��=��.�ځ��&���P��w�
�"�Ob��~A�ֱ1�EZ��G��}X6q����N"� �X%�!�҂;N��
��)�{[����R%y
�}���xy�Z=�ÐFI���\��*�|��Hm�Y-��>y�ٰ��.��7UQ<[	�#����+�*5:�==��(����:����܌Hgw�DǄX��q��h�{��S����s�5�.�(��2��C���q4\�LV��x_���.��祿'_'��,�j��@X#x{֢f��9���&|�Dp�D����
�=��	#�TؒR�?8�=o@X�Nj���gF
Nywb./�'g;l�Ϳ4�"?��~h�g�a�/�q�?V�ݹ:��)'�2dq|u�G;�W�=��`����ϋXW��y��NS%vP$q�\N�,�]8(k?�N��@��H�W�c�*����ҧ����vW@.�]G����U���R��Z���r���51G�i:�&-�ak���¡�hs�G���U��>��=G?�T�h2e�ɳT�Z�H�l���W"�	d����A��7���*����(\i�|���*��D��M�o�	�߇�}]�6p0��	�k��T���kǯ�:'_����lM�K�HBk��y]����"��H,��my)�Y��Y����nC<z5o�8�	#����Q��k���cȿe�?��k�4��$�J�&�6���eʒlW��?=��Q�:���ʁ��Ҷ�G�L3Ɍ���#~i�mZ������-����V�k�>���?c S���]D����O֢TyH�Q��m��f�md\Ş0`7X����54��� R{��t���!W�B81SqZ��arU�����Mx���V9�fb��o^��=��ڮζ�\���ߕ�D6�,���lO��+<*7��@������{^N@�6jޟ:�k�ݟ�,��g<��<�a�$�CڶC�,a�6�A�Ś�4�C���T�"4w@_�@��|��;u���-u�3s�2����ǾLWj0�Y@?���H����	b�U-�G:g,8#ʾB�	����i��Y_͙b�+��4��D���
��3�C0�.&� `�8��[��Z���Hgv>���Vv|�L�v$��}fs��ݖ�[$ƙ8E�,!�0�4�7��r�2ŨlZBL�gd�0�><�\�b���;e����5=�8;*�;�̾�c  �o��P>���|��]�&k����@�/E-v���qzL��G�B�!�Ɓ:$9��J��D�+�����q?k/�s�G%e6>Uw
�����?$��.��;�"��-֓�=�����<G_�̽��.ة?��7H�U�F:���;d����ll�O���Hho�#��*G�XO �`�"�)�