XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��͙Y��p�io�Сe�.����v\N�I2�l��w�%�T	��N ͷ��U��78SDΟS�'A��<�zZ�5X�����+ 1�ѩOYǸ��Y�{I�K/�h����O� ��/���K\����Z���LeEU�0������@�������wv@��yn����Ԓ�`��{������¥Yk7�C?"�a�%��JGO��8�H^1�NN]+9ȣ����
Z��<�V����Q�N�
,J��I��(�IQ���qhNN�4�F�;�R�٥v�ř����p���v�y�����V��OyVN���J�[H���@����N4j�.� ��I�^�I��M)�I=H�泀7�6P�3����Hs����X�$��ZZ2�7i	Wv9�[�6��mrL�(�B�$�/k+7�ߖI<n9��~�1�pd�����T��|D��z��U��O�@�uNa�iJ�5�k?r�+L���^�y[q'�~��
U�\iveq*e�B�~҉K�#�*;U\�׫@,�A�3`O�%]�í��w����_̀�^�:��K}e�"�=�����"���s#����~'�,��E.�
B]C ��vZ���K,g n x�J�n�m���j��W����h������wEA�=��#8H0�U��!A�Zc��*騹2\=�$F��(�-��Z�a���Y�B�{���^=��R�򿉚T/W�	��@��6���%�[pķxW,H�q��W��$"E���翕$XlxVHYEB    a037    1fe0T�rF���rg ��DM/��B+�cq���І�jбPB���A�e��t����R2�t�]��6'sNf�8<���L��-�EK_�b��h��v�|(��nǁ�9�vY�j�6�]x� �-N[v��n��5;X��s��ƫR�aߥ����^�>���Y�l^r~Q���j@H.��͡��Zƾ��z�y�(/s�W4�t�65��9�F��t�M��L���[ �M�.5TT����xW�F`��O���-�E/c��k��Eu>��HZ�϶{��,�sR��;q�9��`̇��wT��8�壱�say���)XLP�/	^K�˫������w!^G}�;T�C�T�+��>(j���&L�(_RPk�:� �OqQ��w)h�WVޫ�41�%~KVoRV����D(��F)4u^��1`���U�k��p0���sQ��J�r z���%I�؃�O~뉳�0@(�獛���0��4Q>����%� �C����H׌�Oi�������c���ʧ4��ţ�E�&C�4�<'�_Z�8<�(�VX�[2=QH'AI;��� x~�p��kv+���?���$*��0;�L�R?j^�Sɭ멞W�Ʊpm�{b��X=�7�e��@[(�� ����^�����
��Ib�!w�4ީ��u�$:��' ^�V���)���^�a)�;��	,E�=a������2��1mvw:���h Qd��f� /��	Z*���M���.F}�-�0=�f��D8����!�E�B�^��Q��c�R�;��a��%��Υ���?���.IM�Uȕ���1W�6��εW�0���p��2ۋ2ҜU-���X��&�5AT��C��(�VL�BI��V;���D��O��@�\�i�7@S'�Z)�Ê-��
MZý�c�ema.�'��^[����e`2�Z���>EUv#Z���������>�XUJS���Ůi�
�N3K?1�_��\Yc��4rZ����"�� ��� �+&뉦W� -�̰1pSް.��Tf���-�L��,.�J/�=�[i�BX�Oc�|�f	^�����N?�ر|㺖q3�*��[�x_����0;�B��1gHIH��s�gb	��$�;���=�]��-�I�@��`g�PO��g��@�'K��MR��[����a0���uv��"��*�U>E��F���Ch�c^<d1Z�0�ْ�ߪ��3	�7����p.Y߲���;Lb�&kv�%w'�ݎ��\t�x�szf0�
�+?7�*��,IE!�S�Fj��C��HR
�R�\e�������^P���3�ୌIa���K���������P�G�a�V(�*���}�pS����u|�`������u�� O+�P<ӈ�t"�پϠ������9oq��M՚���f�j�勻L$�S8���
�UΜ�_��N6����ax���N�&�=�c���%\��&���;�y���ʞ=ф/���~ ۺ���Q�K9K L�G����j�yw�.hD$�%��2O��6�k��K(���]��Z?���l���{�{3�On�S�1f�c�,{
��byq�<<b6#m�n)���x��vB�!�zN̅:�L'	
&o�?�~��,�[��-�'"��i�k߯�t6+��dx'MH��9j��p�����B��Ks/��K)���3p�*��L����+f�SV���y�����C�\Q��gu#��*!lCb[9^�o�ՠ��ſqk�%���z[Q�h@�P)�g�w�HH@��M�R���K}�Q�����d�J�z\UJ�Z�'��o�����M��X����t����F�I߳��4o&��=�em~0��5
����4�Y�te��ƀ{�R��>��N.#)b5ڏR=2o�B�A�zGCk�x���~5��p-�s�ة 'G��<b�F2�z��s=
���˟{���m��y
�vG6!	�h�Fk�O��5�\4s�y�y�O#��Ts����'4�*^
a�[Ƞ�������@�N@�g������{I�Դe���>J� @��.����w�`!`��Q!��iw����B\�Kt]���j@KV"�F���d�|<~n�YJ.4��Ӗ�k�(�`�0<��*4�W�Sp�hX�
Tn��5$h���m�dc�T�д�/�����;�8,�"Vx�B��;ic�߁簵���(��К(A���'����H�i�:疩v=� ��T;����c�u�D�~��,	|L�ҜtS�����F𺓜�Q����+�9h؂�R"*NW�d��E���hߩ��bZ����#(��.HJjKc��cˋ&V����o�y�A�qճ�B`~�������=U���,WH�6N��Iv�l���|)ׇ%�t���S#�گ�cH��B�E����i��Y��m���:��:F>�[�b/W�(r~&����F�j9�8�Ws=O��ż
'ٍB�w�l��k��\z�0m?*���������ub\Yјm;���XU��>�Gn@ �gR����
\�7�0Z�c������.�o��
��j%�V"R�m�!�(�kd�Ad�{j�Ţ��x��@J��MJ�y,��3����D�^Y��J��fR0��2��]5�b}��"�(�СMf��IVy(�m�z"KKL�`�gH]�u�m	:.��P�D�v��u_>���� V6�?!�6;p��f7XS������-�3���
�:웟��}���۱���Y/
q��f,2�p�t����-,��(g
n�!�լ�*=a����G��	� ��ҥ��h�d�)�����_�C�^�a=r�{7����d�ֺ��Cr��J�~�`/"���՚���7���?i���8��FeB�|����2Jqɛp��V�ܹ�`��x ��Q��@�`�	�)vI��ܪ�g���לz���v��H�O���a���&~����V�@�"��2��6#�z�X�X=�X��0#�@do�]��̮Ƅ��jPە!�\ִ�-���Ş5��#�7�śg
��.�eA]�v\��}\zOG�pd&B�����d>�of��Lfv�»��r<�Z�4����.�������Z��:DJ�ߦ�)��.0/Ak�F��z� �F�F�;�H)�-\'��*��Ų�"=�Z*�3ᱹ+��[�0�K�'�
F�n�Oo�"�X���y���rl��nl�S�'vLI�Xj���q�ߪ��2��C`y�i[��XK�p������*i-�����i���f�Ω�s�A�2�qwK*)=?
�vL݇Ȯ�xџGu"4�Ѕ!�\1`n ���g�EЖ?G)Ƿ& ��y翄�M٦���PS���*T	[eX��3{V�|es�O�]z���i�ϛ�{����ho�:98=L�U����	SOr�c#�|�XE���D�Сw4@œ�|.�s�\y�o^"׈5]���a
�'"�m-2��?�q�/��J,��C�ņ#f��v�I7n�g��aO�nf�F��4^�`�q�n��N�tM��`'�6�i;KNkV�����A����N9�c�9�~)��&J�U�5��ە��l~nt���*�@�Xc�8g>��}^q�n�ϊu�B�dYW��ö�z��eW Zr	�Ӽ#Hp��^�c�	��,l#pp�!��sG��Z��h��Er�
�nO�"m�̹o"�#���0ÿQU�o7�I�Y?0�0�"1x�����d���r��n�ؠЂ� O-�Rs@j�\`i�V�E��^���G�6�1t���!s�L�!�vo��Zx�fc�6�E��w����7S��K75cL��E���>�(4�'��u���ثlhs:/BfAOT�~���ř���;�	��n؈�|�Z����Mq-�v%�(��w��׺���rΙ{+�ׅ��la'�\��0�u����p:����ܹ�)�0GkT��-v��C�����a�.�X�u�d1aQl6�_�~F�)yT!�I+I©����9�֝�%��P�"�t7���Ά�_�E��b�P+�u��6����e���M��_�2Ԁ���I+�;�܃:1����_�&k$�����j�k���<�ޘO\�ɇ�dT1"�����E�M�^NH-�B�-ю����α��a�Ū2��j8hEy���j����Q��� �PZ[rN�7�Q�����qo�_1��6Z��ғ�K���%(i��t���O\̌2�7^yM[�B�����ѻHۗo�jyݔ����x���H�d!�ܿ4���j=�:�nj)�"�愾����IL�諫7���ve{���b�+8��A7A�3p� �ʺ��0[
f������2i&���Yd�d��U�~E�e�1�b�z+����ƕλ�D�37q��y�H���Ѭu����-�Ԧ�h��_�W��g���7y�$����/��k�*�	�@|�D&�����r�w@]��sLʢ¶;�M���`�5pC�P_�؎�)_Iw��]J�5U��Ry�^��L� ��`HU�PnX�f��T�V���)�\IQ�2����rW14[-��a��A?��C:�BΎ��u����t�=1��b��)�<Q�/��D藁�\y��C:�jXb
�Q��?a.���4ය�H݊�|ݩ𴇎���v��`�Y��Ў�r���� ������!O63hWɆ%�c�<��ް�,[=�mޚ���!ڽ���\�2��Z x�p<�6��� �j`@<��ЀrV���-��g#G�4hP��M)��2�4�j+Y	y�G�b���:z+4Fs��O���R�MT'L�����)�l��)��(#~�!l���`T���,H�5�B4l%��)�M�����{U>�u>/QZ��@^Kb&g=�F�3s�Sqjt\�4#�E�A>,�~}`��f�o�h�^�]����v8G�o+��6�M�,T�TE �+���ǎ<�h�g�3�x�rZ@$ �ppiX_�,������Ax9���G	���Q���ǡ1�'Yا%i��c����ȧ�Lw��W���q�	{�w�J��{� /��i��&Ȑ̚1-�_o����{��!�1@V�
�9��������sX�A��u��#�z�i�ʮ�X�)}ѝ��0L2��ņ��d�ret�%5K�����$����9��l��WcW��S\�<��%q����e6.�G�S^�g88��W��V~��V�.�I��3����_��s�7ĽVvJJ1}q�?�S�`���F'�0����]�jG��6cԃ8D��d�tZ�0U� ^��N��m�>�z`�����=&���k�	�����[Q
q��چT�����f`��Idݎ���;^�!�@թG�1)cO���@,�](�&'c���0\���F��/@��
i�н�gB������c�|�%�Qb���6\0���|H�%��i4WV���>@" ɡ��
ֻ�*v�Zf)K��j`�52�1H�BȔH��m�������Ns��t8*4��q�BU�/��D"���I���-yV�{KT�d$��O���i�;�[�h=�߰�GA��@��4#T3��ǈ��ղ��4�Y��S��7j�F�;�g�����Mܕ�.`Q�E�s���Kt�t�<	4X߆o�S�7���Z��r־��9K���:��h���0� ʰ�u���.�:����:ډ�J��/�?AҾ�t^����*^@�[�H?o���P��������'ݘ�T@�\�&�d)�a��S�-�o��٪���ʌ�,G:���,8�~��<��Ut�9١�(���@�p�����O���b�yw�V�=m�Mǰ��E��*B;r�	�~��������!m�E�!�a����3A+���1���&"�isu�?�ـ��Z4�b���U&�9aց������;O�؊GΤ�A�T'��u�����|8>k�L�2�4ݚ�d���8�$���F���K�?�ٖ�imuCŬ�Lvt��c���^��M�K�Q^|m��b09�!��נ�/)�
��g�:�b]�����4�/k�!�Dw�,�n�b�]�H��u�Vt7�ps��j%�a��}�_K��E�Q��	�5��Mq[����/9�򗭢��/����3���>`T�T�]�h�kt)�#�:z8�|�(x$��~�/b�!�z����*6�H*��r�6]l���+o$b��c9 �n�@YDV���ճ��}� �Y�\Mm�zF$��_�y݅hq�3�Tݎ�B�$,��CDlB�s����	�M,h6��ȺUy�u���oڈh�������_w�mQ�x�~�D���/`,ld��S�aU�C�J/Z�m�}
3�&z�I�bv8�@��=�^���E�L��t�y��?)�R�q�:�4-����k?>�WPP��`�I����������#;	Z�}��b����ya�Z�A2�/o[�-5�%Ԧ�b	���r%��"6I����V0���6ER RX��GC~�.�ir�[3]��BL�;�,�p�w�~~����S���@�l�"��e>����x��z��2��%~J��Q��`ӳ��"�k������D�wL�F�_y�|�������d«�W�ŷG��9�ǟg1��~U	�V8B;߇�k�Qa7�?�_�C2Y��ۊ��Rsņ����9���t���\���p�s�����q����������ʁ"yA���.¢�>e�h[��[�9O�F|�)<�5b�#��.s�/ǀW��b�q��n���q��������4�[�F�
��q�땨�B�b����1���^�(GٗM����AH�g��S��4f�Ք�Sy�>}���6zJ��d���&�����Sm�O�(���-E�)H��E*�*��0��VJ,��٣N�g�R�n^z�R~Q���O[#�.�4�������q_�W�f�C�U_��d�#�qԠ�-��8J؛Đ�Chb�\m�\(C`�U���Q���!�P��]��s�����n�����Z�#m�S^��n���7�&���[�l�o�#�cC��Źei2V-��ݚ�W{�m��x���5O�sH���)]��а]DXIu��e�03)��s3'4V�\�S�$�R9%/]���R+�x
�td��W�L��>!v������̡X�6�=��f��T�b�h��TWl�N�v?9 �B<W�5jM�w`���#����ed<}���PB�@^�Nq���)�rl�[��)3'���l��.Ƅ���8�4*�I;�c0����G��(�����?`�Y�Z�Ҁ��}��AU��סO &`� U�@5���M�$]�|���&�ي1�!���{�,�LIS�l����75L4;�cZ�m`�e:`�G�/9�"�zx�LOd`-�~ݒ1�7
b8t�xI���E��HʘL��|r��I �-�V4��	@gyV�(��f�}r=�ކa�ke�yx��_�gS�,���c��_ˊ�n�r���_�Q��S`��E�@_�p�?�w�(O��b�g��O�ж��;���t�����~���������sӘ�[���	�̽��M3_��&�K�0�}�o\G)���F
~k��1�vI��Y�<�M�bv9L'���%-C~8����Hf�ֲίFc9n�Qls�Z�[9&3�n�B{��Z�A
��wUW~s	��:�}�ڧSF���M�2��@W�����ҟ��ǒ�>B=':�o�BM7|�u^��+��j4p�JD0Ը��W]��v�l�B�J���`��	:�����%ܫ�Z>������0��]# �(��0/y���ř��[�Ä_����.H����t�{��W�/�̦`[����$�x����6p#+�Z(��A狡6�I���1�W��w�L?�p�!y����J���i�MD~�K;�0	�L^|ʭ�֛���Y?�=���&��cu�����x���5�QPh��SI��G��|�4�HЯ`{�[����� �M�$�ua��K��lC�����f�Vu��o�������q�肗�IWY<��t5���n�/1���8����l���f4�