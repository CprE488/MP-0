XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%QO��D4���)�lsC��%��]�~���ٶ����U)=W��5�@���ݛ ���d{Qp8��_苺�Hev���`���I�X�p�}��������>I�KC]�zc��ϕ(��,D:��j�(�����ˡ�X;�3�B^�D�1��O�g2Ɖ�*!nSEԷ�T��wF:�D�BYh��h@,�����[�i躙]룁{�M���R�P
}9yfU�:o�ͫs�q�F��o���g5�ZwG��f�*y�fdT�k�&*n�U@0On��B�/�Ő"YN},����B�)�#��H|M>O@�;Umtė���t�0��[�  z7`~��S���i�I?���S��Pm�/�k���h���p4@�Z�����Hj���%B�܇����ewz��ULVڋ��F�^储����EO�����|�>�q��4���3��E㺣�΂���7͡���S��]#�,���>Hd�ӌ�1c ���C�����@�oD�B����x����+�vU!O��ݥic��+�_]�3���. $�������kfp��?8+`����9{}���^�Iٮ��w�*`�k<��m\���Z~��8`��������w,C��2���*4#m���;���c���-$����y��`e���mn7H}��|	��ܣ�
Kn=k$���TF9FN��[�"�Hz`,)�陶;!�p�C���-�iC��g���McEH�i��7�*���-`�)�o��>����\�XlxVHYEB    6346    1790Md��h��>	#���DZ}������%Ϟ�%�1��1��O�W_��oR3�#aq_ �d���>L�-(��M:;��Pm�c�~4��̜�����*Pխ�U�1R���(j�����&�.�J�%��m��o�
H����v2��7"�>�[��
��2�Ξo��,��P�	Y�r��Pڽ1\����'�� c"wZ岑�, Rb��فʕl�Ğ�e�u�?�*����p��OL��Y���.���/���ǿ���Ǩ\����̶�m1�S:���"�C�,l���R`a
(#��0k{(vk��Э\B%�������D�4��`����_�k�4Ik~�:;��=��@�_��X�D�'����ˁ=f��i6qU4��$� u�&ٮ}I���~���\�g�ٚ�NU59�2.��(�K�-������ _H~^p	L(HӪD�/��6	o���I��
���_<�;s��@$�D�$�-� ���?���HJ�O�,h<�V$R���1����~ۦ��������U?kV���˦XsDFhkf�:@d"Ay
m���Z1�9����	���V���Y/�!��:�谑;X��
�9�!Nr��w�N��h�0Y&��N�������~���@��f�����=������Y��$�(�s��D��V�'��S�$fJ����Ny����ѕɰ�S�W���¡F�y�lr�C�-Ewg�r�y�p��� ���[�+�Y����T�����,I@��8�p�|^�6�Peo����=���6NI�$!���M#��A�rW�>�Vфy���lL=���� �	�qs|�?#L=�j�Rw2�3w@G�Q;�`@�jp".��W��ml�l#4cu��*��i�IF?�lV������$�(f�[*�4�D�{x*���Gc���$]09Ѽ'��l�G9�fA����(;�g4[t�a��n�{�*�?<�bHҸz�̐|n����1/�XjgO��9VfPhRx15R����_D���m�K��;ҁ�,�_e^:5���@؋mSӕ���R�ѿ�Y��� ��%pX� �a��6�a�N���
vQ�D ���h��-H��bpz��Wȵ����y�+��_��:%,�m�ʏ�V�P�<�N�'��f3#�r����~$a�mS�M�
��
py�0T���$��Z�0�[����b�S@rt�2&�lK3F"nTe�/��Y�F�R��k��g��g-6̕�v��๥T,�܄�ѸŶ�n73bCƆ��*O��ȷH��<�,8�@�	0�m̬�h�#5�7C4t��W�}��*������]���a��Q L�gx��'6�FW�_����e�B����$?"u��\SD��j7|H�( � T�J`������rXW��£%�:(�	-Cr�.Ŭ�/�HM�"��4���L�Mƃ�Һ`��� �]�/p��^hry\�.]}D����}p��E���`�ߎm?T�U�(��	�������SZ,��ɏk3|�S}�:�D�(B񗮐��kV�n���&E�R��6j%�9�Pw���9�f�v6�x�*R���J}E��Rp|�D۹���f���>uG%B���MTO��ΏeE��[�6�0-dֳ2Q/Q;�2$�X�����N9W�R?O�A�F��h����M�˄�
g�i�q�q�M�8ʬ��
�۳��*��~~G�
�6иfyh6������ ���|��l���oI��x����D2w�;��Ю#�o^�iQ��p?!�e*��&����\�^9����Ũ�O2�#@>-k�K(ut�I
� �^�����f	��C
�=Bx�M�����5&p��NIU�"^���=���V��'N �u�?rԮ'�D6����{��_�M������!�.n�de��Wm�#���[�)�DC1Y%ַ���JŰO���oc{dR��H74�{9ZM�/���p>|�ɴ]����y�.����OH!9�d�ͻ��d�'g	'��a?�œ�,kH�����rp�l`����:��&.��B�by}�<D}�,��M�t��;����}���e���B�=xڞB�F��М���7G���l;g;J��k�/�3�-�Αy�Gg�g>�����]�o�T/F���Ma$��c{�nQh�J�ݩ~�IK:��(P	��j�=�k�/eV呸S�I#��Zd�n�M/jw��m+C֍Y�T�E��1�`�=-:�9���!�"�F�~?sh������ק_��t+c+sQ ka/IcI�����=��M����t����@�Y��Z�@�����	ds%�CF���7�wQ2�m]KI�Ta��>N+=w���1�G�<��ʹ4�9LaP j�����Wa����/G�&K��10��zޏ�D�r��'fcKl@><�_�HO3�%v.w*�y�c��O��0�s�#Xmo��[V����A��$��{���D}�w�;�qQ֛RB�%�5sx֞���G���Fzi-���t����S���5�r�{�R`*���ng?Z9:�1�K��\�Z�O����V��/�*�[�f]~����)��G�Ɇa�vL��� +jEJum�p���R���\��������;�U�9�4rf���5�����6t1�-Ư��m�(��� ��õ��ǅcE�sXj/�"���h-c���}��Ð���63|�AJ?�;�N�
���b\���f3�B��Z9;�$^�`��1�y�aא�=ou0ñ+��{�	=������3!J<Dx-��sGH��e�C����(g�M�������	ַg��O��]�m�j̤;	��5�F`��vrH�	j�U�c� ��j-�z7ӦIC��9Q/N��Rj��lo��2/ݽΒ9յ�p���#{��Unc|�8��UÌ�3#����E�f���ʢ��{����P(ة_&��H~=�P��'t`ݏQ�f�TϏ�h�L:�Z�ʂ�$����ӧ��g��C��Oh�ߚ���Q�>QKJz��b���6v�t�����#}�G*xt%��f��S�I0^��P�*�.��K�_=�|Ѷ��?�@�S#o�D���� 5�H�����?�Y̋��h��}�������/����5�烙��(�F�m���T�4+F^wBSo��?�Ƈ�_��\R5nC�S\Č�r�t$�$�|�T��C��+���m_>(cZ�hu{��C�}��)�	0{�	{�ў��#�/��"h�l��r�Q�@|��s,w���-�.]�_�0�a�p�����7� ����)��c1�aQ�Jf3�j}n/��B7"��:|��{�2 Κ�_Y[ۊ`�����)�`�+Ꟶ���壈ѧ2}N�~���&�J����/�IIk��0�2a�rv3�A��|e7����9�	<8�h�h����t7l��Q���_|�ص��h���g,g
�������;��]���}�3:f�$!�(�RщF2� 7��5�J�sh#AۮO>Z���eQ���r��0^�l���O �����@�:�y�O.;�f k��ʃ�8�z�.ͷ}$�w�G�G'�wo�II�"��GP���L~��67�<��z���哽��rR�R%RĈћ�]�����B���Z{ �I��(�+ϣ�m�P#>btb|�e��O!��	�Oyr�� \~c�A�u����Q8t��Q����]��J������� ��M?q�G\� �:�L�Ȗ�|�W��=`pi�ii�k�y���h��~�19��&t�0��X�t:ZX�_�����0;M�Xx��OO� M1"b�CH����]>PS-B`Uz�.��Ym��l����|b],���NXə��D����Ş�IV��Mq#��f9-u��C�i^�������#1M���=Lq]�L$>s��QbG�F&_����I{�l���?�D� =�D�De��
�o�"\H���;�tK+%�d��R��8���KvJ!��Q�T���	��*�q���A׷�|V'�%����^�����O�(_Ozj��m )����9�Y
�W3�?`��F�аs݆M�߁KV�����F�b�>�\lc^i5ol?��/�_��2}ayb��ou@��.A����[���/�gR)&��`y&S��{�2�٬��Rːn|X�aӇ���-��T��}/��%(S|�㰉��t3��0�ɭO��߅�?Z��pG𫄧管�������A��_�0�.3��7�@�K���l'��l�=�ц9l#���g<¥v�����c�:�w&�h�"Q*���ʣ[	�`d�~M��"��ǃ.�WT�Y�Oz7ˌķ��ҚK�gO>����nN�Ga������~7�.*6$2��R�����IE�'�6���;Pjƕ1-x�����ݐ�6�K�q|�Awg*���x���N�9Tߺ���V.s{} ·zۨk�.�WV�:������_�Ƭ�u[ �Llh����V _�Ks�L;�WC"z��IM�7����%�fy������+�O5�?�"4!)�hM�e~^$��V�Y�tJ����Qw�C�І�`T��+�K_���o�����0�ι���D-X_/�ZӽtF��t&�l�c���&{�3��:��)Fo�YmU�lLЊ�Vks��4����|P�r
Ȉ��1�{b1
�%u�Ό �N{/K��"gp��k�ɝ��.�R��S}�%�FtuNb9�QwY�Z2�ܐ����5��Ȟη�F�,�������L�b������s��ZD��#'���T!���)�Ü
��J�e�*�����z�#�E$�o��{ÆN�k���Qn�M�/�I����Z�Q���S�μՃ	���� �ѨKо����C]��/ۧ5�j��zq"�fs41�B�fu��~����X��#0��;��8
}^�
A�����}@3yQ�^��&X�<��L������i���4���x���ti�0R�D�� ��ˇ`�7�����U�b�� MDh0�L��m�.LI��h��D�l,�ۡ����X�}�4�"�5�	id6�Wȶ��V���a�w�����l0(���]"�}�N�7W?ݩ�*�D����e�2߄
ʬa@u���H�SRU88���|
8R��$��eΡ����~{U&�T,r\���(D"��� �n�T��} �c�c��%m�ɜ�,r��V-�q�;�;�!��l#a����ϴTv�Y!�K��HQ>������1A�dT1��kYhĉ���0f�= X�bU�=Μ��fD��'�e�y�5'2�/ʀ�Q�.�-�N��z�ۃ����8������*
�o��+��XS�l�n�	gީ!�O2=�Jp�$��6���i�};��DO}���W:t n�	XT�rQ��E���:c�{���ȃVx�_�:{gJ�s̴^zڜ�!n�^qy�كQ�ŖBr`���B��0sCEH"�K�˱����Pς�rkY��Ӡo���%`��s�|���t~j�o��,�� �GͬZC�����[�7�p��ݻLA������'�!g�1�����o���i���s�:j�GG!B�#�wZ���a�e�������0�-u��E�\Ǖ:��w|k��w���Ȭ�a�\�bL�y�U��,��jl�&���U��]��^�Ƌ=�P�y��&��IU�Dy���}����#}T,P5��*:9?r��M4��j�O�U�E�Zs��^$�V�o�4I�8}�)�@�L٭���P9zC���[�OT�\ұ?{,##<(���f�Cb;�ǔaR�bhI]�|������2xD�y�12_���?aڧ"��>��B��� ��K{�)��#�V2��_��G�C��V�fZ:����n��w~O9S\=��Q����ۻ���|r'�,)��r�X ����x-��g{\��b��T�:�N>��b癀Af+