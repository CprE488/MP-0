XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/�+�3��;\��c@`�mŉX�{��z�b�]g1O����Ҧtó��-��D� !r-×�-Rs����el��u�l�� �;�yA���b��,�)�xc�;R��7�x�f��C�{WQ9����c/ ��W~36J*#F�}���=@o���r�d��������T͜�g���D[J~�E؇|��R)��)�uW��[�ѫ%P��2���������@�
>�I����pZ��렗C��R���-��඿'�!ޭ�G(�-d^Bk{9��|ZK+��P%� b*�:B��[vL7t^�:'g*V�`���	�G	ݢH�a�+�`i�l�a�N�ȃ_��rMqk�ᨅ-�4��� 0����:��q���j��P��
���J|��ŵ�V��~Q����p�W몍.A��"�e׷ǉ�Q2�eThʊH
�B�	 �<���+�t�O:�`<y�#���q[7~��a���)|�o�T��,�	+� �Ɓ�*��n�� �o!����YR�7X_PK%�T��_2V�z&�)&��-�ڣ����vM m�<9{��W4�ge�S�9+]⇂hY���UCG��"�,i �,�]3�:(f�5��fE�᫳;�/Ýq������ =���������l3�s4̹�v�Ԗ]�q�a�JJ����V���t����0j��Ls`�_ȶp�+\(�J��Ll�����
)�*/(,��{�\3��F�T٨�$�o���R�Z�_��.0��;�Q�9ݢ�/C����\XlxVHYEB    fa00    2040 >����7�G�;��i�E2�dz�x�-���1%Y�! ��,�=0��G��D�9��p9��w<�j�I���Ai� ����ֈT�)���f�79��P���i<$��ʱ����v��"�X�0k�lH1i����\���ҿv��i�jh}�-,2��t�Q$Fѝ*׭N��/���d��6T3���I�B	��I|�Xpcup0Gn)W�Ԑɾ��<��U}��T���		���w����$N�c������MK'�S�IX����p�`�K0�Y��(A���j��7�3LX���g���޲�/�
��S�+BA���~���Q�&�9��O>�H��K����EL5��sr��Tup�l`���p�q�nB�ǆ;�HS�Z ~�:��=&�����H�����n�Ȗ��A1��^R��er��I�#�^�(���u$����l:w����2��"5y�q�IL]5�qN���˕SeM�4kΝ&��q��=�mK9�ci�2qU�_�ڵ"���I涙m�V���1���(ޛΚ�J��"��~��^�����r���p�@M���%" d�b��tz]
 �l�$������Q���Oj\��붼���"}YՎ>@@{�T�y�5]�U7/n�p�/y�o!���nolJ��2���Vr3��{�u�zu�-̀=�ݟ(��/��El�eD�)R�>������ݞm�~�ʀ�q8�i/\������n����
��J�fh�U|_XE�ε����ҽ�7�'��6����CZ����66�L%'��]F�(��B�|����Б<a�z�^7�]�����g�g�:_����������SH>&�f�'�X�#�	`���O����=��I��(�ŕj�+`�������*�W~��y*`���#�}v�ym<�Hwj�r���E��h K��?-ٴr~``O.k��{��e`���k�V��pǕ���FS�:��O3C�ߎ(�r��������<�\�$]�5��8M�z�7I�Ӥ��R�
J@���٧8���1��C@^NN���0p�:���N�n[+a6��pv�����3j��{{��z��
���֎���o
���b����ܬ(,h
+�^�Wp8�]qL�A����L���ěk��I��T�A�^L�#R7M�����=��p�`�y��?u$e�i.�<w	�д�x
��N��lt" ��Ԛ��;O$��l���R5�n��ߖ�����l�]���Li�z�^��X�R խ&w˾j��9h/��̖2i�� `�vrP��¾d1�-�7��n�u�]2!@��c� �w��6hR�
��r��2$���yE�"~x�]T��Kc  �?��3�	L�8t��-n)ek��RL���ȝ5H~�-8�����l���\�W�qS��y�t��=;1T2D��+�`Z.!Xj���g��+���p�RdU��ZT-��d���5�}k�Y����N$��&+j����AiIR��Z�Υ�k���Y|HP��5�x���ܙPS'��'�*��}a��H�@� ��&�̧�fS?'Po�C�@��}��6��l �_�ϴ�9��b����!<��Z�������G�v̄�'��e_�/rb�S[�.Oq�k�+!���8���=8�-E`��mL_;��6PAګ�b4E�5o��`��碆t�D�Y�]�ǵ���M�GS��{B��@��xzmp��s�3-5�/���Լ�+����KW�V���3���C3Rۿ(���e9ҬJ��= ���&L�w4���+�ښ�]c�
e��H�Mg5b�� �V4�[_W�*� �	:�_q���4|�O*�|B��`��eN���2��S�U����Z�ɓ�L�$�z�e�[f���H�rt��A�@�N��6
���Nh����.��V+�c:�Q|�9個����]��|��������T̄���m$��ڿH7�TU�(��D�"`��AA[��H|tȿ w����|�D�M76V�Sd��a"9��WZ�$�\���[8�V�����T��Z:�}e[�$�G��S�v1�r  2��۴���o�\1.��������!��=�\�ְerW���\__ӸuH.�a��C�SӇ�,���Df��Z�cX�h�1|2ʨ�Z�����b��ѣ�#z`1���&��B�q]j��f���6iS
�1m�Wс�=p�j,/���~�D�m+��x���]����oZ���:�9�̶��R��(&Kþ���;Ɵ�	�M*�j=�I�����ed���E�S�6�q���%(�_]T!2`�"ٯ���DE GuӍ/y^�
m��3I�[>�F�qo�bYh��xH�0���.H�e�b4})
;n�(��;�K	�ώ{�<���Ǐ��S�4�Jn�����7v�[�;���Y*)�#'T���گ$4nhh+c��F��� x�����x�#V��8rޟ/�hsW��[Ӝ��xඒ0�+�b*�ۢ�C	���"[X���Z��,�M���{�_{š�4s�T��Dҳ�K��D̵w�R)[�;��ڕ�7�~>� ���F���lS$5ͨwI��n����)�N����W��މIQ����l*�MEXkʓ�#P�B�>~bW��L(D;V�H�SF�f!*���R�S�v[���5�j9N�������j[��8���0G ;eO�0�Um(��mz �A�$�}Ύ9�����ª��k�ɉ����Da��:�W?,��qH�#ݬJ><kj|�nD3�h,��<^J�\���^�����hoZ��_��Fp�L�({,�}妆v���9(U��E\dؘ�Jc*#�䪟�a�9�.g:��=dC&@�)Mﶒ4F����D��eb~s4�|�Lu���;l��8젰��꯻�D�E�D��B�i��K멲H���������ȴ���Oc�Qr�yǖ�W}��w$W`]��'
�=_H��l[l)�p����L����`�x��	 4-p]������>:�$<�_�T�C'��OB�7��Gl�B��jK�� 8�Z~�����H�Ky�Ϡ>��uH��#��m�u�x�E�T�-��]AI�Y5vf�_L�[�K�>CI�L��k�Hs�$�����4.����p�PP�����#(k�β6 �3���U7�]h����#���O9�S  QlC�SEV3����'yYME�n�l�D�I���H �Mn��"�Hn���'zZ!T�=��S�Y�������^dѴ���3�"M9���.�%�davOKo:��˟�g�����&У~N�f\q��ݸ��Bn��W$�oܯgҚ� ��ŉy���;�D�����l͕�}�VyF��3���2,�75�W�d���&�	����	^�'Ӹ�Y�o���ܲ=ٜ�<k.W�@	����U�?���N���];�ɏ�fH^�D�k�B�ȏ��r���J��SF�1D��c5�a�*�Ds���N.��=u/���r�,���lX�&�q2E����M�ms��S�=�k�����&���M�$7Gy�]��]��7h׈��g�E�����}�I� 3���K߱VҞ�}Y\~�*0щe�Y6��y���ϐJ��i����ڂ���ZE��"¶��A(Y�|��5I/lZ]	�{Ⲡ}&K7���c����:l@�'��Iڠ�_����v���~jA(�=T#-�@�S����X|-S6ǚt�]�za~��2��Eٕo��4���U�����{ad�$�n�U�QNk�ͼ��6��VP`,��Sϣi�m[��b��O�Ok�f��|A�mF{P���&���<�jQO|1�O��^>м���1�(n�ر�	�.�@s�~Rn�l}�D�\�C�.&���㮨��L�	��K���L-#q�(ֆ(xʪ;�qѶ�1Eal:����=n�U�}�6�b�H�����w/�-�V����N���5	�%��ϹV�0RO��`���N���yo���LMѪ�v��8�S�"-%�!k���qL�!��=�gJ5����,Gg���,cX���x��6l�0^�H��"#��O.=��=��I�C/�����]�^CQ�<��K��}�/^����ŵ��\�д{o����!6YP�V�p�:g3�O��;��#���p�P��/is?P��h�t&��v@>5�Y���B��2Z���w�C�C:���ơ�bJK��@hSl��^�ٱ=����Ru������1�I^8�D���.Y;�����F��>ưr51��9=l�-d,u�(���@J�^ű`e��ֿG&+ȟ��'�,�S�t���r�n�x�����x(��ݻ�'cp��Kڞog���v�Vw�P+��$�1�
��[�x�}��HB䙝�';�
I���T�g�����!��%l�����T��1�C�
a/�=�k�Y�N��#km�i�H�i��	��^W�l���,j�2�M���^�Xs`���E����Lz�,^~֖�_��)�SQ��Mw	� �������>[��`�1��2���Ӈ�u����Y%�]�Mjx�_��;
�-�=AJw�EY��Y��;���Fp���sS���Pnx(�d�Nv�A������n�"eE�f��(e��������S=[(�Rg��O�L�ǀc2s[�W�g��J�X7V7>�_ǝ;u.��LdX���Tgb*�u=�:��Iq�#�`�S);�g��#f|cG_=�m�u�,]�d�*��b�k�4��_��b�/G �k��4";vV/!���}n~3ym��D��g�$
�zA��U�z�P3wV��� ���R�^�{ǜ1я�3�19�Jw^�8��r}�����W�z�4��e�R0����+Y@Ju�I9�������S6�q[y/�#q���$�芞`��ϳ��W��T�:�|Õ6)<X�&6D��=�g6ǽ��_��E��\��Ia��m�l����M��^�����>��Y̶�e���`X�2�=���}	Č�_4ʕ+⟊tA)�A� �U���	X�>���a�P��J�g��h�	��H'����ʘF0j��|E�����EP����s�c���k1�Z�NL�-"���׌��_B��t��9Up�\�̡l+�8+0	TS�ik��<; &ײژ�H�^~t�"Lo�\�ȏ�"���'^�=QV;�~��Ď��1�eb�kVT2y���;k�t��-�->H�3�`��l0�j �?1rD�Ɂq�PWF��Hp?k��Vjר��g������NJ�g'j1ls;2�k�o[���	�ɴ��Z�Gi:���G߉��_��r�}�+���� ��}����[�+�� �#6d/�����ϓ��wҜ�,o��4�  ٍ�,q�j�����PJ��B��b��3�b:I?\�
pd�f0s��}��R>�95�������P�(0�<�Ŕ�,钧���M5cEli���U��n����ϧ���պ��+����*�� 0�sh��f��ܞKj$7#��Rg��i^�=�R�F�"^�x!��Oɷ'��=�ZÄ�u MXք$���~���@f��?X��H�6�J��Rk��2����.����E�Ь��'q�j�E�L�-��o�+���D��PY��7���ͅ���,�t�m�@3�䔠%b��p��V���#T\;�F�gr�����Z�w���q����{�����06����[l�>s2����:�5�8Xf��h0���U���yl)ZTߤV U5c��@��y�'��,���$��:��4���&�eq��Wx�r�d�wU��rx0z��̃TGT�7`�3�Ƀ�X��d�؄hwU���0�M���n
7�gX�
c��1�u�[�(�T��,|�}t�\�P\��M864�@��#Z�q|)��'\�˸x���@������/�bIb�5o!L%��b��p������3��C�#E�Hx�lw�_YF��=�v^����%��<�q��(���Z �B���G�B���P����Ȋk,�F���w�c���Ob_p��Y�Dä����?z�E�&mZ�k𱹬k�_BM���;+��U-ЋD���ѕݕ��7�Ƥ�����#j��욍4��^��F�O���r�|��Jm����Y-'eݾO,d�ӫ� $0ԓ�7��;"rNp�KioM�7Ð�����#7���� O'�g�tu��|w-C�y5�ٺR:ʚn4K=���X��,�k�Ա�$�EG�˃T٬���J�������*�]Z�h ��Q��[u�۝�&i����-�sd�Ą�8Ƅ�Jș�������>	���UѠ�c�s��uI�u�8)/ڕ�LG8�@r�õALT��O{����=��>+�ڞbs�bsRI���=P>�g$����pd��<Y+�g�q�G#�R�n�򺽬�2{���ۭi��V�)����l�I�df�U<"�R��f�=Éjʸo�!X��S6~�(�$�ȫ6�N���ض764���h,O��7b��!�i��L��\�!lz	yݵ "{zL�~Œ/�d+e����}cc/W����h�|0�V�i=6+*��d��=�g�o��G�3��0�6=£s>E=��_J�z!���"��wG+6o.E'F����_�6�N���j�@�47��\EQxo���&�|�s���ǜ� Z0>7r�H,l#@@�H}�ڎ����;+�|܉���+�@���˖+��5�c�喃ɿ�E��F���N�<d�� �\����{�K�����Y�^��w�>�ޡ��}#���Pf�
|5�p	�i��jU;�nDqQ��×�p�������b��ykFr}��<3���\ӏF:&�]�í��p~g��Mxa��K�nƫD��n.Y.�/U�e��Y	O��.ِ͔6�SU�:5ENb4D`:����Tl]�`��D��qJA��,��cAe�������L1fvp�O������Y�^��|c�L+5�$K���zޙ�ߗ�2#i�Q������[cQ��l���������p�Ư�y�[�޳@I�ǏDE\���F�)�$�٭!��ה�".#D\m�**橲�i��<�U^&u��a�f��7���,8fE��mV�6�,E���T��Y���bR�8����\����.H�u����s��]��]��	h!�*м���L��*��]���|h��)�����^w�JzT++�
���-w-���
-^S��s@�M�3 ����a[dg�� ǿw;�k�E�+xKc��-�Ӈk�J�E]_c��e|���@���a�������=ʳ[���L��<t9XdFH\�A�y8�\��
FW�����E� -��z%=��+Ȯ���K�/���g��л��֎���K�I|���q�|rn���- 1�̤om{����ZP�u�i�T!�����ډ�Y6,���)�� �ƃ[&^֪:�
��-�˭u���[��]�|q�$&��a������`ɘ���Ř��0C�ӻ��J<y�����/��=@ȟ�@�)���MW��bD��f,��ITUw�,��*�7��Z�)ܧ}C����J��d=9H�si�y�5ާs���FN�U
��GK,*	��s]���4��:�����b#�,"v/_t9�/���_���ۅy���9vAo�F�|�X����LjQ~�����90%Ð3�򯐥3`8/ԥ�0WvV��AdL��{=oDW��T�2�^1�LU`VC_������ �s��o��i��=��Em�-���������X�o% NP;����\|$����K�5����ib��e�0_s�̓Ɲq�ߜ�{�~�ͨ���D��y���pM+�#[c�YV�־5��o��6��m#ײg6o��[tF1@�*4m���ܛ��6Mf ��;%��Bw�ܔ�<���X�WX�:AA��?�urA�Ҫm�
�%Ā�h�\��򪉽�j]�n]���{�N�	Ԝ��Q�|��8?4V���@RҌ �9v�2����8�}Fg��y�R���Ըrd�������к�3\����PE3ƴYf���X�i��f���]k6V+�(<#l�Pm5��#*����pP���6�Y{U�S,��P�[,"y�
��6G ��l	��}��&�2'�طp)�&&F?�
D�q�XlxVHYEB    4f62     b50T�!�ǯ&cg���|�9V3MM&�nO/(�����R�T�����ަ�NXF��V=�&P��%pE%s��*������q��/N������u6WM��Hko��B��j$-�]jV�|��b�[��V�w�%�z>+��׽�&�U��%F�F����/_�h��-��3���_`�v�\=��a�}X�Գх�P@EhI]�'�_�����B	�7��ڪ;�y���*~l��/&3��oc؈���)�-$ֻ���!X����|%K��:�x,��J�V{L� �K~T_r�k��`nLO�����E�K�0���&ü�u��;�& Yz���/Z����5���r��U�*v�N2�����
ě��GepDV�>���M��pt ����=5-@0�}���k�ؓa��g:����?J��o+�W�,��Sw�Hx�g �?N�W���6�ܙ�tܒ�_��V�w���j�Dľ8W�q�	�����5�fJ�.�^��k-�9�.eQl& <�/&%W�G#����SG|��Bnb��.�1K��z�܀su,˒A�?�m��d���$�K2Y�ѡ���	���I������x�x@�k�R4�/4M8��(��2Xw拲'2dL��'R��\e�=��0kaCQ�y��d��..j��n��c�lB��Th�?�JbB�I�1P0��a>GB/n�-��v�šwo�����2�z���~B��S�.���w?��$���|��v	ˈŕ��!z�Eʊ�*���!=� �������Hɨx�p�fw�����!]-��^�V�o��3S���z
)����̕����?l� ���!!���}m�Sn�Z�fe<����v��[K���GB��q�=���M������URk��P�,jt�{,���� �=m�� �W|N,�ͅ��M��t��`�a�,�3��R�w6��4fy�>ʌ��N�X��&?2�b��A΃cث���h�ý-����-1��\�]E�[c�p�֑��~.���>#�h���P%nB6ˏj5�8X@y�,Y��ll��*������
��s`�Â�;'5a��d�&X�;������\���zW���A�F�ϒ9���^;n;�7E& '��gqV��l��-�-;�������t���WL������-��ؠ��j�lUPм	����~�vb�m��R�\m��Y>��wuH��1��I�ݞ����q������ѢBQmx��6�N�K=Ӻm�w>�oV"��2�aR!�N^v�|�Y���_�9NG�C=�Ԡ�BY�O�1_�pPMq��ٯW"��V��$��ɘ��܏��F�D�,�U���s�2@�*���q"�:��4���;,�g��\��\:� 1���� p	xj@)�D��)�Q~�i��֐(4�[�
��avݳ�ò��*DY�����x�ִ�f� �Wx�)G�1:�@�ʤ}mBF����\��AY���@g�b��3ή�cJB+�8�^��&�O"Yy@{�PQ�	�a[�tJ-V�1֓���F�=�7i���1��!���v��dJh����r����	t����R���<�H�ddl|w����3�I
&�U-{�Q��M�QD��]E)X�Ή�c�:�e�~�Tf3L����:,���������8�J����j��ʣAJh݂��v�ӍF�
��ΈqD�z���6zG �zM����չ�<*���6i���_�aI�����7�ޑ��K6���I�T�\ѝ?�5�B�8@����s��[��#���[�u=��^���ԓ1��1�t@n<�W��14�PCbb�i�����G8�[�g���Q�uL�E�|���U��_�9l4�ˤ�0R,��o��BR9QM�&�/�Z�pdo{h�Q�4���'%^!f7��S+j��e��x|�+ߩ���D��W9k"?mΰ^�WΑ�)!��x��g(`1`y��m�逶.,*"�n�E	L���>-$�Y����<!1$�Eȳ�J���$�Rސa-������p@�?�u�!��-;*j6��P�߽O2��J(��f����}�&�E;,ƏUt�ijlB��uf��=)�/�'��roi0��VӴObT�hV�0i��"z�n3Uw=�鏯]��g����]]��1�BsR��h�Ɇ9]�H��1ĥRkr�W#S{�7B�?�Wϱu�u$���#��f}5��P���p�-� 	���q���(�Yi�F_�[�pT���t��Z��c�L��������E�d�pš���SiM����EUJ�y���	�Ъ�ޮ�V�tà��ѝ2�}?�����j?ʕږ�qO��~>Xw�}V��V�(��=��~_"D�܄A~Z�����D����4��� ��wTe�
ގ�CsqпМ'�N��S}J�X^�8�������wqd4 E�:��p� XQ�'P��)�4�x̻��肆�F�[�������Z#_��[\;\~�`�Z���|��fZ���Ꚓ(��q5F�;TT��,�0j���<������lDb�rE�3�r�<X_�����3�e�xmF���4#�B�x`�H��֛eO�!&|��K�^��Cs*z�6�lf��2֑��i3y�d�kA�g*w�9��Zv��n���!tD���[f*�F���,�	��!TN���y�רۄ柒ia~dVH�; �27��+2��`1��鉦#H���}�ʢ�JB��%q�����x{���4Z�wr�.�ĵбIJ�$�O3��G�9A�*20�Bv$��R�	͠CS�_����⢗�4u�w��f�x�9jB�����x������(���{y���%�ޤ��?�_�,\W��k��;ڳ� t	���_ �l��0���CF���