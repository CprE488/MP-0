XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ʻ\���vVG-�䵏�N�q�+�U���&%�$B�������'�ӎBǱ�(����GO�&t���G*@�� �ۦ�!�T�s&/���/���1�'�|S��.^����j��LG�?�;+������C�y����-X�r�>竴)�͈e9�z����PzD9>��ϝS2�,O��C�C�
�l� ��[���&��vo��p����A�)�;�	#V�����߼k�2����6��-B��\3�𺝯+کd�N��ﰇ�cd��Bb���gd<�U��WW肻�������R�?1�����'�,�f��X�O�='a�X�F�S�8�s���}gҘT*1���e�=�-:m�f����)�V�>�iU��o��Y@��@��,��˽s��K�L�I�Q�^DJ��?�F����#�M<K�͠��gt�����_y�|6y���I�̡�oﲋ�A.��k싆AW�=��d�hO�D[dwޓ
o�fc���!���qҌa����ޅ�:ގMg_�!Y���qi���
���!2�����m�-Ŀ $gi���b��e��R�;"���x}�zu:Bj�Y���:0�����G�weh�tv)������Rm�D�V����9��g�wcJlI6>�9/W�^�3�ʺ�{��^�po�H���فB�"�����W%���y�tӥGwՉ�s�z�'�V���(�;ܼ�cl��K|Z��G=i8sW��'��ѩ~#@�:�L�w�P�/퐲�՛��8�ӎXlxVHYEB    1853     810��)��A�������.�[���o]�B��S�4���ȼs�ݩpJ��BK^9�yL`ڻT�ӆ����`^�W0���;��l]�u����Ҵ��|Di��9����͊����2�˗���P�������K��� OPBA��.Q�xL5?Q�Y��& QRr�rl�ԍ�F�~�IΎi4ȳ���[\�_3M�?�	�M�%ֵj%����Tխ�p�KEy�Ú���\ȧh#Y�@�U��;��3��z8�>B�����+נ3��O�ӖQ��We\.�M�,�AL@�S1�2le]ͳ�d�gH�����&���ւ�:p>o�T�AϹ�ⴴ�(ä��d�1��[әgf'����'I�7�],�T���3�7ͤV9'�|3��Ƃ{�A���-J�(�d-��P�m������SVSC�|̚Հ^Ϲ�:9w_:�g_�i+�RV�pе�\�ZnI�c>(}����ҕ)��X�������
F�I0CU=Ƽ>��׆��ď5cjy�(�����X�A�p��*e�����KZ�MNp�b<���0R>��l�aL���׈s����3k1%{�h�]���/1�g�H�/��0�#0�R���s���s�Wc��(�6�C�2藛X %�z:�C��ˈ��;3
�O_��tz�Vi��-/6-|��	�Uo���͏B���m�؞����V�;I��x�3�b�_C9�$Q���3*�渃���q�ɲ�z}w}��n�u��,��p�c�7Ӕ^�b���,cLD�g�5wD?oGBt�/Í���/J%O*��Pv_�4�bb'L7�1�9��*�tf�ݯf�=�Be�x�w�X�h����1�w>����e���T	����&D���H�s�c�87-�Je��8:�I����c�ErM�OIv����aZ�X�;کh"p0���A�i)�v`k+�t�	ɹ��F�3Ӝ�$ܙ���(Lqz��<��IY�����0�^7�*���S�L�>�j[2eA�o��%��>w>��ç߶;E�7�oI�x��*@젃"��Y���ǰ4Ų�Pp�o��B炛�_'�H��f,��0%^S����S�[~�<�A�FLM�	\���ni۬�k�����nt��\]U3����]e�dK��i�߰����SWM�k�I��a\I��u.?5Kiu�y��1�/�|�HU���̨��H�Y��A2n솂�ރ�!B��� f(���}nf�4e���v� ԡ��jR�/Z{�%�`���(%�}��L�̮��\Y}_�D4I��`a{�U��������!s"0����(���xt���H�; ?J�����n�3%�c=�NzY��5c��BU��`�d��aB3��vT�����3	'�i*�~��*���u��>��}���$���]��A�Rs֑0�w�8O�
���@Hʄ��p���'��08�ܭ����F2��4������)�,c}u^�/����t�xM��H��tnf������ɳ?7d���^�J�5�4��%��0��Ϙ��O�@߻A~<&�U4�MDR��;1�g�tv�����qQ��(�V�.f��
O'��g��A+���^k��5���J���B�K>E�ڀA`ߖO�M��8����z`�[��iՅ>z��}l�XE�ɶ�b��d8�؁2�� {X�w�[�t�Ц�dJO3s߆��:��u�gc��S�n��Ze"�=�}	��^72�k�r�_G�h"�`�A��p���m,t�� �y�h`��'b�: /~2{�CV?nS��������V��?v_S�(;����ٚ��iT�Er��/3��ʄngey
�r+R`6E�FZ������< ��sv KL�pտ���次{N{Wt;�3\����p��1��`�O�u� �U���	^�%�Ћ���c�7{5����v~p�R��p�|�pn�̐��j����_��[a2��A"Z3���+{~�αl�J�����=�$�S�����������e�v(��u��>1�,�����D
[ן��WҮ