XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}�[��XUAh�$�� H��x������x/'3Uc�ʏ������^A;�h&A���q��m��cK S%>A�"�Q1M�׮W�xa�
��O��v5mB�[�3�Tu5��9Ii��-�^����PF ��ÒT��s��k�պL��XToy�^[���mm��{��T�ݚed��|\�>������v�"�S����snn�K	�tAiIŹQ.�TyJg��Ͱ�&,�RY�*Ї�:�'��=��^�6;����}d�~go�G>��C�\���jW�w:�mV�?(���u�݆�ɛIh�O�&zi�O$޹�C�s��u�T�fLlҎ��-�8�[��ú�~Ix ��*¨�iX�3�??4��V܄�{(J��晢a��2��<�i-���g��m8���8b�P>�s4�a��O��I�ig�Zs���=���X�����`����q��>d��*��)��F��7k0����\Y�>��f切a��e�Gg]5�#N�_��g�?�j~)Z��q�>h�r�wn��!��Eh�|tǖlIe��DN�a��4T��+n.o6(�m�7��m�?[��쾌�H�x�3[UL�]��N��l�ʦs�3R�ps��[��{;9��%X��[Mz>�V�߾�q���~����-�w�)?I�
��Z_t��H2=���C�,j���1���Ue��_�5ٟ�i޷d�ur�/7�z��j��)�B���:�I�ӧ|�����:ߗ����/S�ޘ<�j&�� %��XlxVHYEB    a037    1fe01x�����A���ʄ�c�)j*:���ز�y�ς�X��!5���Zƣ��.�[V8��O�Y^�b�#�u��@��+����O+�����t�(�x���K`=�{�]q�hF$��[`�qX��,>��H�����U���K��sg��8��Wo����MX������'*9��X2/�8I��%��)U��cTT�텷 銤�.�Q�מs�1'ϴ��C"���c3���(��y�!���0P��RjB�@t&��v�2����'���ol,�+�����#�C:j���O�
���� �ִJ����i��J^]�ts�@?�S����M�KW��=�����;�GbK$��N,x� $L�!��t��:�A��O���ې E���R�֓<D���2��+���b�>w����5v��J��X"ʅӚ 71R�C�y.��,1;7�}����S+���-�Ƚ�Է�e1��NͦM&��e��%a~�\��4���^�L� �ԭ��C�d���EP�!D�Ũҡ�=R��;�X�(��z�����|[]�UX_�b~m!�7�g�@���Ǐ�ѧ��d����g4Ȍ"��w��m�Қ�	o\�,!�:���@C�������:7P�w�u�+j���D���M;�scc��
L�R�H���zfcA�GԼ�~;�o��:��P:�՝,�Q[��b�ľ6��'���3#	�D	������C��)�_ ����y�(��7�+���"��q5��D�j�(F���<���5�I:`��	�^�N�YĂk�����&�)�OxܘLk�q�����X�P~�[�:DB�(H�>���$1I_+��v1��d*'��Y6�J�+�}t��e�4d�!�+Ѿ��oB˖n�9{���ڻ�<n�f)`[䖹�w<�����r��G����8/�#l��sh�
������93'p:`�H�w�t�*\��Jn��m��X!X����j%ҿQGh�C��/=gǙ�,f}���O^��Q��o�AX��d �[\+��$�2/��*ׂ��ls	�TY��<,�;�O.M��K�WEa5 �X�)��Vo��F�q�U�#O2���@�2��m�O''g�L��>�H�����?F�B����U��IU��a>u��¼��l��X��N�E�wSʕj��$���Yy�SI���;� ��ؘ��|$VS���w���q��J{�4��>q�7a-K�s��Qt��( 8a���I�)ࣹ�c4՚ġj)�[�e��$$V)�v�0:�Ӕi4�>Yʼ
<�<��ϟ(��Y"L��Hϋñ)x�+���	�أ<��vhDn�r{\�'d����X��B�U����%�2,�vY ��@�LŽ���q^��@P<��ȡI����ўŁf[ѥ*�0��� z��$S]��?�jykE����M��躘��{	�N�s��$�7 �sUET|5��p��TD�����h
|4����GH�Ľy�iU��X��6Q��}@�[��p�m9��C�Wt����!���4�߫=wv�T0�V��o����p��N$�U��������ɵpĳ&��M�o�i�Q�+M���?��� Z^T��)*��r�7�bg��q�F�V)��BR
��: 6�Q.�MЅ�+b�����v��{ea1�b����@1w����>G �fާԺ���Vaj3w���B�\�@YMX��.�~G$5ߦb)<�� ~Y�9�9uQ�>5;�e�B��x��7�iyp���P���Xi�m�	��o5S'�pc�/í|>�5r�-���.]⹙�L���ҢL�7�-f�NK�e'%�$C�"T���0<z ߉^�m8 ��[����a���0��]�(�UI�)k�Ӆf�˯�!��u�5�/�-.E1gV�=��+��"ɏ�^-�Y��K�^�$d3�*ъ+ �0Nd��Op���)�!|EZ��M�߯�@)�C��1�a�%_����BsF@�s�cF�m�(�P�(=KedW��TӢ%����/�hQ���qU��28��n�N�0��D�9~�o�2��sO�/�CN�v� �h:rM��A���5[��L��!o<Bc{{t	Ե1G�����d�-.���2�@�_�_��;A��+��`g��֙.�#D�>F��H<v	Q�Q�6\��L�+�������;�j�;���c�b\RkǷL��mU��J��G-�]�Yu�"5�z����j�x��8���O�9��(}�Q7e����b��7\ԅ�*�(w��%DV�8��!-Q*/6�&L�:�~
*� -/���+�����9W��3y�k��׍7!�Bր~ i��D�G���7�=Hr�w�|�2D�P�uRw_�Z����0Ꙣ+@�8�v�E�D_�R��6���ɵ���t#}��.�v��n[�QՊy������>��E~X��0�Hn�7ܕ�B)����Zi�Ϳ��A��G�\�i��GjZ%��n���E��܁-b�y��j����Y5�~�f0��g�]` /�����2ܠ�MI8F�Φ"g/O�#��s׏v\v[`��@H�ݟ̌�C����gP]i1��U���د��&�#qQ��.�̝�A�и^�0�����Z��%k��r�3��I���*%�p�̷C��@g�@uz;K��|ݛ�������td���5�[wu��5�/M��1��~̂H̖A��2���l��F���A՛x.iY�B��jjFk74�]�&^�F�x!wƨ��M��;a?�}�#Kv���G�X?�Jj��VR&�r(��a�}�p��=	�Zh�C�;���s�<�;���i/.|��́��z�n\�-P��$�q<4 8/��9()�i@���"�`�h�[�~����i"�U��d����;�h/w�B��@du.���d�Hh"�B�r�`�䞇�\���p[ڛ��rbnq��Q��F!�?�N�Tm4��wʊ��+����vn���������U��+��yb��#�ʽ��G�Y��"o$z&0�Ns��%�uG���wc!�&�_���/�n��	<�d莨t�2��h�R�A��^�.r[Aq�X���(��}�p^�(��_����ā�ũ��i7g`�X��!�D��n�^�u�Fs������
�lۉo�z]�����P��/:�J��w�O����j&��!�B�:|�0�!Κ�E�}Ǧ�g��������V�Q3L����f��%+�h��J�3Q m/�A�sL6�v�Q����=�����.	'ȍ}��:3?[2}�⸲8�;?�� Ws^"zޛ|�r�ک	�N#��Db��Ր�����p���n��e�z,�D���>T�e�e�n�h�2c���\�!�1�_�BM��x�䧂�I��RƬ���]�e�̵<��	��4�,����B/�[����l��"G�����׻���O�Rt� /�H�ϥ��*��(k���驌P͖���M̱���^~��<-As�՜)$��q��Ԝ,�G�p����\$�J�-
b�< �{�H�+�W���(O
"=[�ӊ���^�t_N����\iB<��>�WB����ȱ�����hJ���7Įq�Aؽu�<o9����ӑ��v�܍��.G�ܿ�\������Э�ī~��M����HRsr����c�X�k�h@����8�!�֥�?qH�[ݡ��Ъ#Ic�f��@ƞ�}d�������E�8E1���N�=�-֜(�v�L赥~���vrw��jc~��� ��c��
)0���&�i/��2dN��,?E)m=KDg7r���t���t����\P���`��e�sq�y0�8"�ɰ����Ī�=�ᆙRQغm3���B,57�c��vx��W�E�x�vxtc �3_YQe�ܤ�R��w2b7�?[�U���	��!#O���m?��΋R�3n�!�*p*T)ޘQ^��r���#:S%����^_N���<x�i���J��f�/�%����0l�p��M���L@�w����!H3����V�A�����GOo��Z ����ܜ{y���ڷT#,ځ�A_���IɿPgWq1Z������>��|���ֺ�%iS�$�c�ыU����~�Nۈ��6g�N�h�w���/�����w����yT��	k��u#��:�űQL��)���_n/l��A�߭_��*�%F����A?�h�*4��c6鞡� �V�i ��*Щ������~��\�����EP'�G7�N9ٴH�!�ΞYo�0=���v��:�g_�! �Ũ���7��Z���3|��*�D,k�l(�<<o��0jӧ���ݿs�5:3B16��,3�N�).9!�S
[���+>�-U�� �o�7.��i r�ȟ�|L��&
��z�v�9�@TS���o�M?��e����:�1gͲ�N���ug�_b���e����D3%���V�X�,=�`��rc=��9l\V�ߜ�L����B�i8��/Z���i��d����Y���>Ҭ���5KG��zQ�p�V�ͥM4dL�!�����l[4Ψ�#U�TSqx�����+��2]]�7<p5 e#�����\�\8�z�@q�&��u��V��D»KKX.��z���c��UJ�+Sq߷�en�x�����S�fT75�kq)i��U$�q^l�[C�����ns�~�)�N�b:��n�nKTH
|3�lๅ�c]TD1���h#��d�#�����M���3�	ҽd�:��I^���Ա)Kl76.{d^||L.}�����=3��q�Y&�Y��!^7<�V~zy��?0ː��gǧm�l:d.h�����j��`�;��;��0�\��H��qC�!��E@��8��ү��]�򎎿mGF!��;R_#���$|ܴ ��so:�?����.�!5[�p�����D��C����M;���q��W��b�d��{`Ǩ�V㣽Cl��<���F��im�Mg�h��9�)	�|
ʫ��ha��]�^��sT0�9����|]��K/n3�؝���8����%"Ө���%��ݷ샋�#�K߱�'�C�&ǹ��ܱU1��s`��HҒ`��B�*r�ލ!E5a�t+\�@"=k*$Ϻ�������fBY���C�M�sx��� )9u'#����
�K"|�y_T{[
��3qdNmZ��gҍOd��UM��V�y��y7��#2�p�a���.�j��6�_4Z��V��ܢ�V����UI�`R������'π�Ӿt�a8��#�`I~�ڢ���~T��R`���H��	��Z�sGɈ�4��\<ؕ�t��H���d�1�.H3�2p:�)���`�r�-OF�����3����^uQ����;����Y�q�O�ޗ�_U���Р"+:j�w�L�H��!<�i��O�>������ƝP��ʡ1���ww�J�؉��X���mn.4�,ʴ� �#YyÔ"�:������;��̀���`�ݗ���R�a�2u#��ދ���������b�F���J�AV�-��O¢�D�X���{?���BP��"�>�y���B�����K�K��(cT	q��C�dg�V໊7i��L
�W ҡ��*76�����Ϟ
�buAr��9˫�c����:�:m�H'<FH��U�;V ��{W�o� �ٝe�0�g�g]L��I�h�DZ�D��ʶ�3s_�l�b�l�T��d�t`�$�:.˅�,,QW�,���_�RA�'���I��iR��ג�w�,�b��������r�9U�+��[=��f���=�-^s��(��TL�0ujh�CO��a��8nOF����ǚ[p�-=X[	��,!��C�£���������ђ�/9����R��6��Ӑ0FΘW����t)��E&٤j@G۩����g��m�diF1���+���;�p �.E����Umd�&��t[��`�AW�Ra}t��]��2��5�����p��n����n�Ƭ1�!�w�U�� ����Tr$�����F5=��e��$���nj���O+"��6^���ȩoPuV��E,�J��pXL�rG-��~	'dMa:$��.��@��8�4	O�1ɔ�<�mP�D=y�;?R�УZ<��&ъ��41��G�ME�.R�"X��/�9�V9�0�'���V8Q�fe��0"�rx\��y�fV���x��Lvy�s�dVV�dAȾ��������^��+��}�{��K���F�a��n��_/X����=z��ց���R���_�ᄆM��r/M���݇���	E���QY��ڇ"zc1�gc�[��D�KXr�ӡ��Gzze��zU�u��zw$`#�7�̒V���*z~�y�?� l��D�@7�M.�Pltz�)�A��n���4(��j�����*`�7�Z"峪�.��Ć���M�����e�\�+Y]��3���ΰ�z��/H����k��aq�c� ����;�?}��]>�M��B���}!�9�}A���H��JE��x>U`�������)���GHY�͇5�7�T����g�d�����ӡ���##(;D��G�ٜ�sW�.��v:��2 )>}WF���T�4��k�\Oikȱ�8b���O'�_�u�L�}DM��x�:��U�i�'���9��7��H�fLq�:5�n=:+}G���? �'�~��Yz��ոbԶ0��R�D�����M(��0�M�Us����E�r����lW�4b��b��/��6V��Q�qyM��W#r�x �?���47V�w"�g���ڣR%R���G�}�n9!тe�l�5�0�y���r��G�'�g�cq~CX�?���7�?iZ�т�o�k.��Bǥc{ۛӐ?�r��S���� �"�T(ǜ�ߝ����(�2���%�5�NWO�̔�����Җ=���"�������g9aݒ��Ee�4/�1qF��-IX(C���`�?�}�����@��\f�/x��$l�:,������G�r ���l>�MĴ|�J��k*�Dlx�s�E�Y}\bM�W0|�De�+!:�W}��m:9��@���{�6sDN%��SAT�e*����J 0{a��ۗxX��W���� �`�(gJ7�0�w�k^�E$*��	
�����w[���oyO��\G�ɟD>�p}n��WC�HnK��s[S}nGKG����x�B�k����+�a5�A���<����[�AU�, \�?�L�K.�t��E%%�#�m����c@sFMo���`���c&}M���Db��Ć�'��%A��p��".��p�> I}-�Ē�f�K�D�B��^�ǡ�T�.g�n3���	�G5"�LK��s+�2�y�X�mV�F��:oK�� �m�#��N|
s�߇�
��t)�8>�eoQN��&34<#A~��~��T���jXԍ�g��'�݉J&'$}R��r��O���v7�����<WJƫ|���a-� |���b���Ԍ����2f��~�S,�-�Ȣӟ��V�<���g�_�{�u4gdϖYE���Lv��4�[r��r�)����D���Qz��)�detY'J���b���Ķ2��C�׊�{�ī"f(k�����;���x�����i��{����B�!����Kؒ�`����@�h����Z�P�8��@��?�P��M,q��e|�3�0��Y<[ĩ���-j�J+�|��l��qS"�'�Q���a8�H}�U�C��%q#t�_!�}��ѣY��hD��}F(�'����k*�pR�f��`9�kp�[?C'�YvsO*�y���~��&��I:�n��o��Mk���GA�K�Sm/S�Mv�8bgd�	��q� ���iO��^�BQTb�̴B_5�;��P�R�5�gZ����f�?i�VZ�Q/-���F:U%o*wL�CO��~�%�S�����[��"����IxJ`��� vս��ţ�i8.�Mv�FK�F�%���"�J�uI�e& �G8��Vo�M��s�����2u�'�e6X��=