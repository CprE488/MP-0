XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{}Y{���9PU�A�8�j�B �Û#����	B� ��}D�\�o�����E���f#��I���;x
\��V��nM-L��]��O��9�Etqx���X��5��&t(�w �|2(�{E��h��)�`��jA�~�ڐ���a���d��'��9����^z�������w	H�����wlE�8��<e�8��˽}�~x6��Fl��S�A�Rp-'Bw���A��b��h�)cx��cqM4�5t�8��I5�8d�ߜ�k^���	Rv&i36Ռ2V-�y������خU����)�z�ĵ)�M��{��H� �q���|+v��n��X�~�_�	�Y]R��!c�8<��x����7��lJ�-��E"�2}yX3�[�,���m���Ű�G��_�O�JZ}0�M�N�O�?��k��!�s��m !�:ɦ{
�cVy�#)`���Xy/�P�.n;i��ý,_�;+���G���[�G�������S3]wѹ�̿{��ݳ��4*� ���3�x緂ɭ���� 21��d7����y�3@���o�1�{lw��X)G��a�7�8�H���|E�12�n��9)�0���"q/�0.�Ư��N����P�!�V!W��gP$�^D-���ް�U�N?�]��a�)�,�c��@	�Xڡm���,��hx	�ũ�i}��(׭�Tu�_^�o0��+�K�:]���*p	 .лO9�H�,M6�F��������kŅ�#1�XlxVHYEB    fa00    20400]ߜoAIEUF��dPO�hkkɔ >�H&Ɔ���[o�%<��R��i�|�@O[�l�6��Y�j~4���.�¦�(����h��d��������6�_Y�L�;�Î�5���Q9�J(y?E	f۠:B!E�+�'�Rp��Y��oW���H ���P� �3�-�6� I���K&��R-����i�h�q�NY�W��IK�����0��v�+p�,�ȀI��}WJ�Dh�f:����q�e��'���푥��7,���*\TB(�}3Kd�a����������i�Zo�4�L~�U!hn��;`����
0`�L�)zؕu �'@�H�����|(�@_y1��dXx��В����U�� Wd�8�2 �]�J�����K�i�`���*�3x{V�r.�n�2�FmKZ<c0��Z5��x�a��A~�����>@���j`v���m�6�&�����Lj�ƒ&��4��Q>շ߼�8�J��h�@�8���|��%hDy�U��P^�݁Ppa�m�����+��ikA����6�C�R�h����c��;q[���Tؑx�MG ����q�	'MYB�����Я�|Zc6��	�������BP0�mٍ�A�w||��*Ŝ��{��]kܒQ�GQE���bT������v�	ݒ^�b��^�k�Y��B*��Ɖ�J2 &3�K��.R�UC$���`HrȰ|i�~'����¶(Tі`�h�g�`U���"�� 1��f;4�G	�TX7�Fݻ��<��*d.�Όş�[�X�����$� �&�4�k�d���j�x�IѮۯm�9�#g�i�K�g ��FN#����߲��t����������`i���؂��?�Sӈ������og�U��������
I����7�87�5g�����o6�B�u� �'�?����[�v�ѧ�*��˟*]AF\w.�>���];t;�)�5i�����V]��j�`��D��r7��ɟj�������5�7��2�%E7������Enp��a�
���<yz׿�Qݤ����g�����s��R�,@L�h�]dT���'���m�݅Ӭ�|���]޸K��*ͱ�A;�L�L�3W�0��Ԡw6e��`��cI@��M��ͬ�(�O,H�����E�LWhƈ�}+�\�gǓ��?������A9g��xU�7�/��a�/�� ��N>���42�M0��
WF�z_�W�D�S��@�=��k��?|��*��#k�y
g�+?XBR��C���9���w�8���B)�r	����nԋk�^�=�rjۊ�����un�%58F
�f�Bu�dD�>)s$D�s��+����S	�d+m�8lR=�tO�B��_7�=��� ��	�]�����,�PA��.�;��m���nb�U�Yi��9�8���R�mP9Xۗ��3�.�є�J�P�zb��{�U�q������2_�'�; .tkf�O��7ɒ �ck$nd��i�c����n�9�&kU��yG~���r1�����T�����r2h���w>�e-𱑅��w=�@e�>��,�9X)@���Bq��\]�X�vy-B�F�ea�@Ҁ���2���	���跹Ք�ZS��� eĔrL.��5�g�ҫ3��^S@��<�k�@����B���1���IM��Z�G��@s�\u�d��FP\��͍�j!7�.=�S�V��d�ь	��v�I��G�	�;^�tl�����'����1�Y	\|�����f[���H�T6���^{��2�@+؛oƓ:�XW<rr�م�7g��X~v��PmV�^<��{�C]���,8�}����~���x�#l笮�p;��R����t��U,�����j�ظ�s�N?F�P҂x�q�H�b��Cg�j�%�7�*WCss�Gj��]���yC�_f/�M��h��k�7zi��_��H��:2b����6?|�]"������@��\b͔F��ߐ��Xa�a�4�ta��Is��B��s
1�l�t�%h�9�����O۴��n��Մ����Gt�����By{�C=����)�1��dT�^���z��Q�[�o�Z6&��2ӫ�v��D�U�¶�'Ą4튊���҃�/j�e;�Nm�e_�(�>�p��AJ�+�Z�����=�z�����CC[� �|I%V;�v���FS�x\`;"�c�V���1&�\33�R��n��6y1�ַ�ۅ*�"�R�Cx7)o	��`�`?��HX��1.�tu@7��K%.�C�����Q����K�����ׄwgK7�[���-R��o���O��������Sn!@��:�b0;'��n��a��d��ߌn��E_�۔�;�E� _\��.�.�W�:�)j =^n3�}�h�w�}2xXR����H��mV}M��nu}�U_������أPI�y�N��N��FЃt��y }쳹\�QC絿A��j�Edz�}�����
��4�0���W�����^��%��Y����%:�-o���p0֬�V��Z���'�^�qӢ�Ȍ��*�u5��U��*ST9�: 3�NA�x��&I���agR���ڃ�U�6ŕ !,G}d���h	L�R�T@C,��h�ʻ�|��?��ۨ�ݖ�R'�W�+�7ȉI9�i� 1� ��l��ԧ��Q#U�>�&�V���=�0���rW��r�ɶy����}���b뀪Tp���G�D��N���r*v���|�`dfĕ�5�R�L#�s��n�����G8��ɀ\��|DT��=$q<?�b^��&7	RI�aXd0��ڊ��Zx$3�Vg�^���^zhO��/BdJimY��GF�[M�x��}��D����>�/s��7M��
�d��=�����Ixӫ���^ q��9u���B�#��}�;Ϲ2�.c7Ht\����u������yZ�{���&�8r��iOrwfAi��L<
�RŮyCd��@g<����(���`:SY���;w�Ms��IQ�� a&�ʄ�7d��:.�K���Z�"O�3��ʏ�؆��w&`�374+o����~{�L�.�0~{����0i�� 1>�CG�:*p����$�&V� � !�x1��g+����LX�1�Q��7=�	=azL�O��}{#���'���e�L����	�����"��'�R�#J�	�JP�#-@��?ָ�<C�C��e+V�{-��^�cQ'e��Tإ&��L���Ufz���JO��Or}����I^m�g5�6[������)t�3�/�ˮ����+ޭJ�Mk��^ON���7mס?�3h��}6�CE���t��ȇuS�w{��}SK@����@���ܰ��e�̫l�����5{�����ܪ��v���	m;��T�������yN�bn(��[�0�:�4�����a�ѣڂ�?�S62�܁*+d�e����9^r-w`����&5�H2·()ӭ���IR@R$yk�V����M����YK���u�Ϥ��U��\�s��~�C8��)��`�*;���2�k�i�Y%e$�hB$�­��
�q�fZեx�N��Z�-/#��f�OZ�;A��lx�'�56�v1��-uւ
:xD��l�����}X}�V܋A!�x����K����Q ���2:X❚��)rc��8���	��Ү��A�-���tZ���D��A��YV��V�qO�'�G�sl�M�Q\��u��[�� m��6W Mo�����iiǀM3��[0Ҹ6�.�
��E����i��aǗ�*p��97�8��Fز��eT@1��Թ�1 Lb��,� �ڷY{��"���۸�=|fKJc��H��W�9�&ZRA<X􊬄͒V0��}����o�m�H�uTܯe����#�^�8�Q��l�샌�pB��U��i�y��-�N�=!IM�#6��{��<i�F�Q��� �-��䬫^1�gNF�{,�2�z�Y�A�-�y���q{�D���Wǧ�[ڼ1~��$-A�kܨc�ϳ�c��j�r�-cE@�K�O�og Eݼ>o戜w���� ���:%�JN4��;Y�j��S>9���X�q�89S*�����vG框���B+7�&��G3\���7�]�Y%����D��Q�m�����.CV��Rr�{�e=R!g�<I�t�b]O�a*��OI�!EIvT"P�������b5LM4]i���;#a���H��~�b�ͧ��1�g�墂��7x��T����Ɇ�n�b^	�ն�ô�/q�y(����	gBf��UEp���+� �e�� lU���i�ޏ#��)��[�DN+v݂9re�"V���[r��d��eLK�k�/�_��������J�@eJ,�t�xKP�<�0�5�,6�Dl�A� puX�(5�q2�Q�m��q�#�	�%�>��]@��V"h�m�+��p2���ye�V�q��	��Ш;��=oPy)&��j�����'u1 �&�j}�KG�Ǹ�c.���� ���K�/�+�i?��ֈ�~MG)��W|���u�hF�2�jP�e�r~_�7�D%٬ŉTZ������4�j@!b��c�;�%,��yG�?Xn\���'AH��:x���sw��}�vO�Y�.�a��1W�vi�vG�t�u���+Th��B�t�v�p���nN3�^�M��V��tvX"�*�����s�Y���M�c�Ɲ?S���atK�<�0��0���~�Ԕ9���^ �k�O� 8)L�����'A��zJ�T��QƕL�衸A�y*�,[��W�L;�0.�5~�*z�W��j�괺���U���.�����,�J����%������ͱ�o�/�aH<)�=�#�B%]1����F����ڛ�U��k���e�Dα�����lp������X&� �tק�����·d3������O�������PfA
y���@iPckw/��ċn��i��:�p�Lb�ȣ�� $t�����Z����懤�ѺU�պ߮-̞��G��l��"�(���.�F�jd��m�����J��hv�m/���j�=��Y��J��IR�q3I"o[�(�'�B2B�ֱD��><ƺj�h�8�n�9��RğIA�qc^�������>�h����w9M���Z�kM筅Q=��w�4ᔯb����K>s�~M�bK�[�F�)jbŪ��*����ui�)�������P�|�S_�6m[���� >�TDt��|�vߚI'!��.QV��C<z��1���*#A�Kξxނ��3¡�E�9�8}���si�����B���yٟ�8�V�í�p�];s6�IU|)��*�!���R�	��������N7H.�1�����-NB��/C��F�t�0)��y��ʶ�V�
 p��@*� /G�+ʃ f���DK|5`�g����%�q�Lg��L�"u�!���_�p�v(�WP�ids��+�ߗw'�T%���ѿ����%cU����s��KC@i�g˲iE���=��'>V�b����GGS ��wӭ9��i����e��`��̧W�;�vY�#�u"gxT.���Q.��f���$)+6��]Z��e��tuM�B����nR�A[&���_+�WY��%3�X0b�o�'J3J
l)v���,�_�n���Nj)T��Ӈ�`�6h̼<x�.-J��N�_�4~_>΂�t�f;\�1���)SΚ��*�K +�/h�}�(7"��S�&�uC6
3Ύ k"47�?�I��Cx�7m+*����M!�{'�?����b�ލ��%^lEW/ҭ���IR�_�`bPo�g���G�{"��.fZ���6Ľ �;�-	���������o�G  ����#���ԝ,*�69�����p�"C�p �~�F���:W�(cbh|*Ñ�����M!����ƌ{H�H㈞��&�h�W$��ر�P�|�y%n�����g ĚKN������ErH��&g�����V��D}�G���h�ũ.��'Α{��[�����կ++�M�۟�_`q"DY+d oeֶ0�J�|7����.DR���뽫���-����R�r��W��2��C�ڏ5�uf>܎��IЋ�F�� �+d��M�$
/>wP���9�H��V7���S�+�(>�	� K4,f+� �ި�oU?EҸ�4js���Vz�Z�0��_���\TW��8l��,f4�M�&���3Yю�;k�oF�r�%"^t+�L����+�ޭ�f����P�.��E\� �p�d�;��]M$�/Z��?G}�j��5������m��ۆ4��A,�m��ܺp *������<�Y��nȈ�R�+V�D6���0�8�3�P���e�P��߀$�6��d%�.�oN���5�W���qǜm��*�m4,g'�Z �G.Q,FC��,Hs�U��?�b7n���M���%8�!,��ܬ�V��U���(�cX�6;������E�^1�kj�ߎ�}@����r���T,j����ƀ)�Z�R.K��!�J4 m� ݨ�[�C�
�[v��h�(0�sF��3!}
˕����.�C�Pj�@� d3U�]06�:ʏ*��ꃴS�4U�}��:��3�r�f���/Y��ڀ�a�U�n@ P�����M�)�R�3y�˚k���~=�.�y�{�0��k#���N�K�����(N3���y�=�W�D���E:���pz4�Mv����.�������'\6��~Y���Mt;:	���~$�o��xF�����y_p~,Wqƞ���#Yg���
�%ә�ϑ���Ś�|��;:ҩ]v�t{l��`]Z��w��Q�e���Cd�#3�]H������l�D�ܷ\���xa+��s�e�+y=�!�;f]>}5WK?�H�A�H���I����S|�\AjK�D�o� ��MGW��-���aa|j!ugmR�����q���,��.t �v	R��U=/���6 +a���d*�]8�F�����"�p`z�*%���Ί/:܄�6��)?�0���M{�bm���P8�Q������������|AQ��L3u�H~s.CV�������s��G�xX�w_ff��1R�<�����6���D]�wK���}Yn2��ʽjg�{e�˵ƥv���!	��]`�����h]���s_�5��&�Mwf���M�.�
oHY��b.�h�~U���LK\��Q׈7�[^�)<�#;G��r�9#��h)D8��״��NN U�8W� n]�Q��ĵ��K �`g��W�����?Skݦf�0�_��X*���S���b�6Cg^aj�]n��@A��"Q�JP�fVOm�#�A	y���^���L�!�Ubn%�Aӣ'X����뚠Q}��!�X��M�]R�pD)�@Opz�ب+k�宲�rn���������Q�	�w/��m��g<��緈���n�#�q��C��c\0֏HN"�&������<~z��,S!+u�7fmt)K�攝6h�dIx����D_��UA�誚��U��{j5��+���<#Wt8At��+��w�������K�Y��:��{�H�c�L��|��`7���+>
�B�Z�bl�M���l�aܡDrĄ�π:
����i���g��H�o� �ql���Y�`_��k��b�YoLFy�1F!S|�?(�	2���S��������k !C��S������f)'P*.A]p�yI��)��9Ŀδ�x�H�� ��o���؞y�F��V�#)�\�הFz�9<�Kx��$���೺R��'a����U�~�:�l������H?\{��B7�UZHu�1�|���4h��$�i��$��%>��#��*w	��T��(RbJ��㨛�=��K�����O�g�U�=��0�4gHBnި�����f�lt�.ɡ�/�d����q�\	E� 잲1�-��r&︄��y�t|l'\J���j�/=�,f��~fH��F�_Ś�����0�V��|:3O^�#K������)s�5�������1�*[��8�N17��w�ϲ�C����L;���p�d
>2���Q	�?i]�9(��#Q������������Z�>XlxVHYEB    4f62     b50�>�,����(P'a6�m�zb�n�*��ia���Е��19E�#ft�9͸5�e�L�{�I�:����I��a�o��63�,:X������6�G$���y[� ��D�F �_>��W�n�*�L�������jC��W�A� ʦ')��s���ގL��F�t?e��ew^ �����}VS̃���OutC��Ѝ�M��3�L��n�e��4^"��>��ӂ7"� ���AZ���/ Xr��*�\Mu�l����;��7��=o"�B�����Fe7�L�:[y�6�����"p@��;�`|X?;p����n�u���6�F���2����H��H��֏��#;��w�!�UJTC��1�5�����n��V^N��qO��������/��W��~(�-�ϯ��k	��2y�D��v��6�m\���@/^�;�!���@�����KWr4����6
�p۽<-��Ŏ��;�)�9�h9n�%��%5��J�sJϨ��:��L:k�q���:SI��F8��5�5��j�DY�6[�h�ř�f�p*&��m�9C�#VӖ	��2��?e(1Җ��f�x^�Æ4uhM���I��N���S��x�$ޒ�ە�.+E��#�!ʫ�ºy5���7�<�QX�'��B�;"�'<����Ýi�uJ�¤���ڮ'z���ڧg���-A����3&f��O½�\�a��p��mU�bm]t�)ʉ���x��ɾ��R�k�G_.�e��ao����1;�ސ�,����_�(l��65G5�A9�e]8	�Q�a0�A��m�e^��L�Ԏ�ir�q<��8����:������)�<n��,�{�-?QS�sQeq�����`gݩ�k~��ŰOZ���*/�^ʦ7)t�`��p:���h�p�"uW��w� "��9�>Zk�xAb���q_��"���B{ZB����n��i�Z�/+[�|w�H�&��_��Dp��J��J���h�������6���6(���Qf#f��S���65�W�f��qvu�3�y��'4��k{�)��GGn�R�Q���R�c_4y3Y����Ê��6қߞ�F�m����e?g�J-�@�te��`9	�RɅly>��/*�d�[����`�N�}Γ����7F�hV���l�ѭ�/
���}�iE��Y�`��o�>���q1#h��م�n������ђ[>�L��G\}{��=|�4���=��q|6�t=�4�61��I���Sq�M~���o�1�!���E鯇�DN��}N�wJe���v5�����"p9=��C��߅_?��X�$@Õ��y���A�|�Mψ��P�~&�-M[^Po�A�}���u���3z@�Y���˴�ϥ75kjr�~�u$�{���s��4
��������Ue(���acf����{�;c��W��-J�#�q�A�
R�j��{�����8�Z�FҸ!�N�1�+a]��	��z��88ޫ,��Xm��A�^�����p0 U{���L������� �����F[`�\�.N��z�1�ZKk��J5Q=�ɿ���"����c����Ml�F{��՜!�e)s<i�n��Rݰh�T���	�)q�s�HI1(��k�
#�`���
-�{E��-��Q�](w�x��y2��?���jj{��&J�J�׀�pJxG]_V8�ڮjF��OE�&ȱ�F�H��m�X��Ґ $9��u�U�O������.��U����c$�(��E]�� �,'�����Ym�Z�Y�ĳ�N�qbd�b���[��X��L���D~��Ћ�#�YΡrm�A�b��c�&��Wn�R�������N�A���(�`6K1�2����~{	m�!���t����s*���r )~���T�<�$Y%L�bK�u�H{kp��C�9�%V%�\�"ﺑL&2��Z(���� |;NY*vyk2a\,'�"B�9H�F�b�ױ[$��m�X��0�� (,ƫ�VJZ3A��c%;=Vb���1�I����jA��S<�1�e4Ш����Z�~G�4:9���e�m�A�5��0�z�Q)�~tEa=�G'��wFK��
��r���5�9�!,�E�\Q��F�Z�^4` �xaAn���67�n��s���>��l;��v�ի��������Q+�5��� o~�ݴL�Hc�Ɩ����"K�qTf��ٛU�Qy��������2�'5�sB�>�Y����M��3<M���w��4��f$琡#y�Ĭ���E9u��g[�f�2{0ʊ����ð�%ҍ��=�u`(�8�j��@n�>]��������|��`����d�����L�J�.��w�i4�%k��:D��%��e7�ڏ�;��&�Ո���������-C�ߨ/�oc��LO0l��լ������T��m��tQ.úymUŔ.إ╼��X ~�:��w�5%�U߱���x�l��8�DI���i1ۗ�6Y�� ^l�'$;�������3�lߝ	׾�OE��7!��wN�y8N�����)��?i.ۄGoV�/mQ�8D'Ed|B�?`�CEY��p��n"��\�m��i1���A�ȧ����a�9#1�����e�|pc�6�>��f�֟>2��/	a�C������m�)7�����
��(T�8��:j�V��f���h�Yy)z9�ym�]��/ӭ���Q���aL��Ĳ��Gc�?���>K���_�4/upA�}���V� �F�R�"#�\Wxa���}�]EU�H�Q\�d�
V*9V������J��2"��K���~�J�^���L�t���\�`��ۊ��;�}a��V]�C��z?Q�gvu��o��_0�d�;�^��