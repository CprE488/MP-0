XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l�T[չ�M�.������ڃ���:(ZG�т��������ѧ��2N��eǷj}��uZ���%^��(�:��H���� ��RT�G��~)�UB�2����O(�;-�񫼘/|ed�����˓!>����y���:P*#T~��uW�p��Z��**�TA���>��z�ȧӗ	�a�v"zk� ?�94V��fN���u��͠Z��(�t�w�d���nk�)=Z�!�K=<\)��*0Pқ����Ω�O�yw��O^Hm|����FW������q0� {��M-�^�:�@�v��|���w)PZl+	ۙ� ��W�a}2_WϮsuH);c�L�iL��yTxZ<{2�֮����3�Tf�O�d?�_O��va]���ʃ!,A51n��P�c�iI��X�!*�`x��|;�~p|!�K,\l��1�:]��7�����T��viiL��"9���u��1�^���RZ����40-�4�CLc��OVM��L'i�rQ��<�#0KG������ ���,�Z)^�c߿�T����E7mD���;f�t�J�"�b��W���黅�n#�j�]�_��V��Gt��+$c��[����;�C(F5۴O=�V�x*�B�����k������]Z���zZ�7��/v�Q�~f߉����u��U3�͸^�>��,�&��H-�u�R--�J[<�U'jr(\"�����C��
3S����O�8 4 <��-�^��(}���G�����ZXlxVHYEB     f6d     6f0v�18�ʫ�t���>������&���zmĉlD��'��ʉ�*��f���%f<}=n���G9�ET�i�H�I�$?�S�u��)�lψѨ>D��C��T7�ne&=0��u*����rNL)����n-�PMןG��h�k��E��� ��5|�30�ս���9�F�JJ_b�x���&��-�g�bO��/ض�w��`L�C�O�/֙5�j+:eČKid�g�Y����cs��F�g��hf�GeU�7�C�	:����@�������������������9�����A(��A��H�I�S�w���(G�^���{��gp<1( ��TBZ`Oy��󔘈�Ċ]n��#e%Y��� 
-#)�����{$8����tmK���^^L[�'���)Љ/g��BC+��g���aە{���;��X��ג��B�kQ�մ��qҽZ���BAr-����겙j�GQ�@9D��l�`f$�Q���fU��� P[3���Mq��!ȼ]|b�,�����&�S�V��>�]Jm�0�_d[o���C��A�Ӝ�Q�Q��afSҳ�� .������^���R����ܟ�����{�߫g����h7/� y�{+Z��|�@�fRN���P7������8���}c�7�G@li߈��FzK���*� RA%�+�Ĳ�g�H�$.��[I�� �v��|�b������^N���G����"����2r]v���Pmb�Ŏ6�]�¤�u�=��[}����r�j�~���{�>�(X�JqP�h�INV`IS#Ii���S%GC"�]yഐ�����)�hmQT�A�Wpkyي0yͻ_fS�p�O�8$��a���a)���G�M�}'|5��oG'��^I�N N��m1Q�a��A�:�!��w�y8�wG�f���&E9��V<]��1+�����w����"��� ;�� 0MQ����2ۣ2	�'Q*6�������8�����E���Z0��-����:a�~�f%sj�(��U�Q���g&��	ۃ��//��eU�(yv�p#9*��'���ln&��q;����]oz #�Cx/��i�Pz�4r�ȕ�V9GK���5I��~Y��w���	D��Q%�����{d"
S�"NW����{H��n(��T�eY#���$�+C�Z#���~Z��/���H��X}��W(Ԋ�O�a�$M�$%�>	C�k����
�� �oDT�Z]t���4�#�����Qd���~�N�s͊�Llhop��Z�d>>�ϧ*�����_8_��Ep9�AR�6(��O��=��8S#���|8��z*�%�L?`c� �h̹��)���xq�s+Ƒ�Q2���S�g75��%�_�]տ�1e��� �y�F�h��yB/��ɒØ������a�}$��y�슎�_��+�=a>N	#���3M��O��
�|�HЦ��"ȑ�88SO.F/�׳̋�7��t���ˤ|��J���;��L�YP�6����� �� �x
$J��k��g�蔙R��>	��(~���}�sяl^?�G������=���F����r����N�ep��(,4�Ȱ-���J���J�����Bj�W8�Ӻ E�<x�F7�[�w� +��%�u��+�����%�!'x��x�d���6]�Nn��F�vB���œb5\ӿU7����'�p������Greo��	CO�4�����t0��ˉM�1�nז(v�{䱁�4�h�``���X��,x