XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���q>�I�8�̕7O��B�Er��y���3��3�ߛ-NqK��Z�J��VPa�q;Q���r��Ȋ
$
B��ԟn��bME7<ł4�
u�	y�G� ��Nbɗ��]��"@�P��AL���#�BIz�Z��"!*�l����B�n��\ ��m{����?S��2}�,׭'`;��`����X$��}o��K����j��LtS���¯��
�n왎By�ª˥Vf�9
�=kp��QK�y�'=f�n�� ��P���UK^�9��x��fu��`����k��&7�Eow�q�?�n�r�K�I�=�?O$U�����Mk�+�b*�ݾ�4M�b��hۑ��;��G9=��IL�4tE+���P
A�����[���l�f�d�V��u�k�	��DU�$|L�{�!�;N�4ቒj� �߶�H?��>�Y1���`f��m���W7�L��7�G�,g�a�ܵ�!��|E�lnʟ���55,6�[�N�J_�G�隥�Q����ec�tz����:���׉�B)qa!��Q��k���'<u*g8��D�Ad�%-&d:��I�~}@��!��N�Ə[�2w=H}�1��4-��~4oK!���!��4�����FN�֨�:&��_k�Ս졸�EɢƱ�>� �p˙���B��rC��jտ��P�?�C�w;��<�x�N�i��a{�Л�P<����R�(���s��a'��;��^�����@���^.d��6C���<����AV��#�2��XlxVHYEB    6014    1840��BI^z����=���>�@q�E!�OZ�oBp��,����TQb��et��;�dODN������h�i���YS����� �IG�[oG%�q�6��e�8���e;Yf<���9D�jg�^��]�.���b|�D���{�N� �c9�bp�g�](Ud�ga��A :�zV��Y0i]�Jʑn�I�=B��Y���mu�׻��:I�5M��G�k �]�u�YjB	%�B@�Z���9p����>�4�o����x������="�J� �
u�QmX!<e��@��)�����������XB�Fݐ9i,�#dJE���ﴔ�0S�`�T��#�Ą+Ҿ�H$.p��;�,p��B}cتDDH׀ϸR$)�w��� Bm~���*�sg��&���Xm�iƺDM)�W^��szP���TC׿Ǆ�����\sg茓l���R�F�Hć�a��y6����?-��hS����q׭�Վy� ��jR��0$�9�)Lڞ�k���t����\<v�-Z5&z�����=RCZ�]w�X.����)�6������K�sO����_Q��/ჺK\]�f��Ā:н�G6#�?$D��8ak�hBL��j�Y�w4��!�u���CLC>x�m�yG�����<���|
M���(����1=t՝?C&��>�[�vn�ER�'s���-���g���	��� �B��^ny0c�X	�wH1���	�H5�9Ү�-�Y��t��$n�s/;A"�v`�r����f�r������Ъ]��RmB?կ�2�|��!������Y�d��ܡ��y��m�F����vF�,j�4|V��������F�R�X]�N+�G���m;����@�e��d����O�P�-p�HS���#�O\S�d�ܺ�@]_=!�x:w�n��*�lE=Kn��L�a�&"��,��`�� �zˈO�������n}+t�:���D�����^��O�m�Pf
�C1�l�{��">
]�k$���?�o���=8��.w��N;o��7�w�U�a���k��D���S�yho�ǙZ,��rS:to��l���5Ze��*�ެ]�>��N�|l)1�m�QѺ�tF@Tα�ҭ,>�⟛�}N\ݸ��v��M�cy��֢hXX�1\���E͊d%Sn�:� ӕoA�9����!=m�e��U�D� `�Y�Yϒ�gK���%n��pE��hc��]�ӹJ	���Z�Lʄ �5�~ek��u�o���`I��@t�̗ʯ.� ��xj���L��(�:<��n��D6$�+�ч�:�6���h���,��oB�j�ܑ��e3D=�׫�B@zm`�R�f��iGܼd�֯B#�X��QS�G���M"&"�J��ߏ>~��aa`9��V����DX�L�cE�~t�z�Eg�?��0��ko}����q@T8~ݩ��n�;�&��L��� ����q�M�S���<T�)��H���'}��ᦕH� ���X2ʐ)/�q<1MC�G�@���MQJ������}������"��Y��>����3�)�O@{����"��%��xWvP�����?qM�{~ �����T���բz��Ò3 �b��T}��⎜,���Y��F@�M��v�}��E����^>o��d/u|a�w���Ip��O�`�٤�2��$��,���=��N��E�)(�V#��P��0�u��3x�Q/��V�����y+#�5	ce�H��>!y��僐�^}��mT�^[���J���V��Js�;�]�,�q>"Q�we��h�(���HkK���qJ�YZKZ|��� ��V��CM����������%g��r<�+��:X�~`P�����a؃<*cC�`#�D7��Kζ�nU���]�s��]R<;L��ܙ�Ә�A��L�2��zJ�1Zi��p �Ї��� n�N���D�JZPp���`�e���j]�^#.��d�.�Jx��y�,1r.}�OtL��(d/��(H[��^���r�4���Ea]��Z�#<:�D��n�?�=<�����Ys\r���dd�̙(��ɸ۶�a�+�v@v)��EA�~\ɸ&S��2��/n�o<Z0��kŭ�rbi��=��7P��1������s[7������!�);���<Vt\��P��4
���P��-�2 P��kxѯ P���&U���S,#�\���<�.[��#z5xk9]�Sz�1�����H?�<��'~},mIL�;^��C���R:6�ub�/	֨���0a��/���S޲��@AԘ�L%�2}�� �__�ț�3�2�3aX?$�֪`�X_
����e}�����T���~��gN��(�G�6�� �yf��c�185He�4�KJrb��h�^��vu4��d�gA|׽u�jM(KM&������+ٚX.��ͯ�g^���0��3�>��j�j�I0k��V _�(�*	��F�5�
U��U��x��-bnP�'#��������&NZjl��XݚU���+ʂ$��|�I�����a\�1�xz��Y� � �5��}u�,�>�:^m�"��g_'}5@`>~�w��t�*P�a��]�VKT� o݆�zOIJ�Gϭ���|��|�kfȥ�OCW����*$��� �� ��=���a��� P����Z`�E�
to8I��V�J~PC���9�h�G��x��3�W�2;i����f���t5D"Sib�K��m#��@7&���H��� ��&�`�%E�W�fK�QA$W���w�5���ɉ�d��M�^���������?�$�-� >�۾�z{'d[q��j�4Y;���ːϾ�B-26`L���V�M�	�d��E�k�B�����vclG�Lj�?`?�$buW��(l_��+<�*��e��Cd�4w�S����8�	ܙ�H�ke	�^�wgi�T��Й"��C�kJB������c RK�N,���v.�NSwY/CO�mC�L�Ws��9���Vz�k��F=�@$
��]��.^~�ƚz�C��&��\-��@ ��1�N�&�E�m�n�����N��|*���q:W.߫.5�8̲���_(�}�
�%O��7N�u�Ss.�ן旻�}����O��/�2�4�2��)W�\�9��>���Uz/���kZ��%g�;�|����o���/|y>�P���+��H���h2�����=6:/�c�*(� h���
zs1��whW�h�tM�n�wVMUןB���[y�:�օ���@��.�q,F��ݔ�Z�J �����]�5L�P�� ��|��s��r��t�ު[�_�o�ln�9$g�b�˙��dҡӍ]ܙ��7��� ���qo����T�[J.�}!2Ѯ6Uh�3a{(˵�?�E����U�i�'$e�:ieiM�p����N���F��g)n\-��>( �g��p�s� ��·��}��눏ܢ�~ǖeN�^��&��䋆|�0������',f���췐0�)9k�}�A��K��"+n�<^gr:���������d~ 1N�Cˮ�݌ɿ���kSOt)�@�<��Y��6l�%U���[!����tu�<dG��@c����׶�\���F(6��̋�y¾����������:�,R���}��*�@��8�Y���=ks^��~�����!��4E�����
�j!�6{b��C_��p�Ǡ��ye�`���{��İضs
�P��:�V0�J�̅P.ΰ���@C�Pez�>���!�r�֐Ww�-�V��v��Ws:��
�&>��&�F�֘a>�0�}��!"Sp4��������č��!{�����ICxa$���q�s���S/K���P_�e�N�U����Z4���*t؊�%��c&� d3�����}1��p�����|;�	Z�\�Lp=�������>)�~g�-�A{2�	ؖ�� F���ꍔ���si�]�r���YΊ�6���4��@Qn�*F�q�@���Q�����R�FP�Is/_e�5\E�Z���	��z9���DŎ���>�
s�er�Q0�o1̛��� ,�}�Η��e5�p�0�IF:�h����V�=iڞD���g�/4��)��qC�?.?r�M߻�������,1jj�Q��(�D��pW���u����_�$j&?$1S�⑳*���E)��7F/���� �M���0jJD��݋�N�xx̖;�b��JU��f��(��M�B��Z�7q^K��%�^.�(D��u�!s�QwA�]p��fx�,���2I �>M� y��v��!���O�\�2��1]��'�I�G�֜��@qD\lF�p����5{g��i4��O�lu��s��G�x�I�.���W<�AY��Gî��0G.í����W�V)4@{<��+9��P�YyU�#��P7��wG���Y.������=�u��)��W�S�<Jx(��fT�p
�F5�L�.���Ϊ6; �cK#��c�b���GE�Fk�eo#@�?�mt�/�v�9�e~&)�G?I���Y#�`7^��)6��/��ݦǻ����/3A�V�
>�W�s�R�D��pI�FOD\@�
�]F�&��]���� �	 ���T#�Oاi�4;����K��(H�R�j���{Ul�Ƒ��x�po�a�97~O)A�5�ŮM��"���n,��N�J�i��	~���s)B�2�W��Hx�V0���:IE
ږl`ߜA/�s�jj����1�t�����x�� ��Ȝ�M�\/�Q�'��D�[%�TbYF�	n�{1N�&W���+Mŷ-��������|nJƲ�����"S�o�}Y(�l��"4���1�RE��&�$�$�/��l�R���6}Y��1g[�:�ٵ$���B̟; �L[H��=�Kf��"`������$�����#q�}�ct�2q'��ٙ
��wk4o|����}'ۗ������<����>$$\g���U�OK�̋�]�wW���K�L1t�]���ʘ�v��̈��Q��5�����.���j�hua�AsJHh�{1�s�J��
[����ĦE�\w�+���1Z��1l *�����"]�8)PQ�3���{���L<G�UOA����\si�k� �8�/�F�Q�dLu5�����6_�E(�EY҇��g�V��8?��zo��7��;~��8
 �7S��u����Pോ(n�Mʫ���e�a�.T=bβ.B�G���թN,�b��� `��vs��������_ ����W�"�$�o �Tv��'�l5�"}`���YW2s�< �.�Q��L�ȡ��vt�&�ghG�7���̩����f��#6�.VϢf���E�LC?��v����:d��5!��7�u����vҚ��uO;+X�Y0�vY%N�;���� v��^��ոs��J��zf�q�w^�4�����tX!�^�%�p�xZ�;Е�N��� o[hwW�j��O���;���A��)�ߍ�$�`b�!چ���E��tKP�1��iQ%�p�$�"�%�\�j��kS�U0kЈ���.�)ܱtѺ���k[2�BJ{R�1��ݓj����Uw�w�-�(w��2�,Gwrt�����V�]��z͚
��lf��L���i��h��9p�%#�EA�I����˓t4=� ��r\�vZ���H��?ȷ!�.*=��8�-�z�7G���TW(ٝ|_�|Jq�L�w��Ib���^"eڶ���&\.넶�#��(͍��%��n�福ej������Iu�O@m�e�[� {ٶ���ܫ rr���;}{5rQ96�b�E�iF}��ƌ����e��m�P�A�i3/4��/���Y���@��*Z�x|"�m)o景{���{:��Rƣ�pl��A ���d�`�?ߗ<Ğ��;�f�����w
�������b��f��!��C)AO�����0{��N�q71�,�����^J����!�	9ͷLz�Û���S$A�9�e�w�b|��e�)|<jͻ�`�8q�����u�
v��74�gS&{TS��N��W�d��؉�vx���&�/�)9q|9��Ҫ�{te���[����