XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w�`���"t�ؖ&��n
���>�����^S�c�]��	�x�QSf�ǸVe/�B�u���N0��o�~�`�}��q�_I%��x7%�f-�,p���9�N;�+6�o"�[�fo��!H[�]�l�V�\[�f�\��b|�=O���'}��I��C~��]��]�_0tAu�'#���e�`�E�چਅ1��t$���G�l-�1�<u�o� p^�Boj�kk�?W���l���L� Y�V��D�V7,}�a��E�0��'@6�� �_ۍ�����֊���O�����oL��'E�Lay�bFH�# ���V�HǷ����=��n{��i��-	�=�p��xE����E��?�:%w�dO)hg�Ȯ�F��ԃ��C���@��:�/���\x_�i�ef�o���+Og/VG��I���٫���g2ቾ�����Ϸn��q$�ʞ�p��mҀ��1.�Y纘���/�u�}�ͅ��.��h�! � x]59ҳ�R\ҹ����D�z�.P�}�x������%��+] �Oz��֨{�'��Xt�X�5�Q��-L!YY6�����f���U� ���e#	�I�|�d^[F:+-aq�T��c�Â�UY�d9��:����[S��=�B2�x�V$~.*�g�d������h�_�ѿ7�ֻ)��V��d�Z�.�5LZ�Q�2����G�tsǹ��.r2Hit~P����H�%��HQ���2��I������\x2�rXlxVHYEB    1853     810�]��k*G3>��V����JG}������P:Ș�VVC+��cj���d�\!hH�,}���s�2���ÞW=�@]CH�8\/?�l��q5SuȢδ��r��ȣ/2�|�X�0�G��}Д�*���UB�8eA0��k��Z�0�9�Æ<��:�L�4���+�XdCNO�
=8�����1�Lp��m:���0�;��X+�<�(J��m��9JV'qH��-b��8���������n�+�[Y6��B*��lR�wO�D6����Sj%т�,�7�A�	�+"{�P���-M�:%�I0g��H#�
@u�.�D ?S���� Hg(���	�m,�Ȓ���n�.��rR���+~	�w�Ud�����a��o�y�2�
�C�}o�)�=��a�S(�1~Į?��-�F'J��K�oIB*�Fry����3��.�7�g3�e3��R���%�M�@���h��HH#O���-w���;1��Û�����1J��f�ͅ��p(sD��^���'���Х�uH2��	��uLRj���?���(���Ʈ���%hˠv~��P�����\ΘGq��M���.��I��yh���G�ˠ:t 9&�]�[ �@�1>Bm�}����ف�@���#�����XV���K�w��$Ay�/QS���$ܓd��Rl�oI���[N�p:�6ݟ
���cH� 3���\_�>c0�	���U�e� K�%he�^�o��J�gqԧ���ۑ{V!��qY%l��6��ң�o]�0xx��~M�{6�k�ă��7@d�K�MG/�����e�r����T�*9�v��?�=|R_� ]�eB������/��?�p�:�V�Хt�zq6e��\��zO<�� �Ps ���ֻt�å&��x,�A�4�_�������^�q1��#odlH9��2�}��;ѫV�������Ź+��7�?}���A��/��fMyl�4�s�k4�ESݏ�������Kt�����WfOuU~'~����$5,i��ɂ<;k�u*�YiͻDi��JE��A�h�<��(V��c8�/�w�,���k��8�Ux��?���ɰ�a$�a���ZJs{N��rm}���:@#�@� @ "�����������D�R>�C!����	(�1�3��W��4HߴK��u��iҙ��yt>��ZAK���.ǌG�-{\L�#� b�*F�:����72t�ѐ<�|���-�� ����v4��I��0$D
M�xG�0{.�Ց�VR�'P��[����~^�� g$�إ�z?x!eX�V^L�=�b]@1��cU���{-P�Ԍ9��# o��x*�n�_`�1�?r�31�m����bՉ&Z�F��>����X����"j�8��P�����'>�b��J��cx�;���� O9]r;�1��Y4VE�-�:r[�x�8<ݫ��F�14<�	#R�I	�G	}5�*J_׉̞W�Z�gᓱ�؆�igec��DK��'�g���bM��R�H7���T9��Z)�}��H�P���C[��S��'�)^�>]�5�m@Q��ޞ�7�C^,]zQSփ1�?�0����{����2�7��r��)�w��슷�%e��7�Ht�a	qQY�z�6�>O��n̤�6�h/ߟ�?����-�wA�-�ӝ��������ؾ]E:�ѱյj�T}�nb��	�Ď����Bl+����<��?��˕=�z�z`�G5?��[n1Zl��"�*�5�m��`t^!^M��"yqL;��\k�zqZkJ��m�q�@ԕuи�R��l�<5ڪ�
9"�3C�م�����hP-gh�V�Ǆ���X�k4����.'����Hu�u�6��q�����y�]��0���Q�o��uQK0�L��K��G�L:Ex�B#�r�(�gV\�j��%��(�G�F3�)!>�fG��fp��S����r?*�b�3� ��Ux�6���%��E�c�����!!_�G�k:�5��3)3px?�r8�2��8���G�