XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���k������hJL��zBD��ߔ���c��W`������R��uV}���?'!�̿������"|G��z=�,���&`�XԠCEo[��ǵ�|�b��H�4E�M��"�73�û�u�s򊚿�4X����WjN�ܷ����.��ز�A)X�A9q���6g")M �M��}휋���@��ȯT���{��e(��@,{�����z�_��N�e����&���
	�o�찪�~'p�j��p~^�sѣ	%v0��C�ҩ��HVwYdH�M��X������RI�'�G�'�#_m-��R� ��*[����|A*(�o�D�V#��0Pn���5��t���yx��'Q�U���`n�F��U�i��n$:�a5��P!����ۧ�RM���ץ�g(S�c
��su�7kx��U�a�ɍ8�+�ȇ��Ĺ�Z/�Z����S�?���|@�t2t�7]��c��D�Zm�_�J����ڄNg(��C�=�a�k�<z�_�T����Vb��!���qg�����é�k�N������+��n�2?AE�y��D[�M̪�U=�_��懫�'�	E�'@4.������E����}��zR%άֶͱ0�� X�^��9��"8�&���K�����ٯ��\�u��:� ��`�f�u��"�T&��'ހ���Y�~	N��S/|8٦�+ie���j��݈� B)���i�(����Ǭ���tӛXlxVHYEB    42ae    1110��l~#Xn�)�l~��o�C�"�x%Ū��!4�8"��8��MR�W�"Y�E���=k�G �����`��I�v�����=��ꋰ�ӄH'p�_b�)��W�u��������"�"���
�R{.}����uC\�ș����v�TO~���z�[����Η����X�.ĩy>�U�D��1	�	�(B��@���[\���zD�����S�z�o�j\�4B���.q����h�9���;�j����$Bky�|&Vf@C�C��)��j�a�
����n
@�2�tz[	��Zz�93�]m�nN����0ۄ@Ƒ�|��c�㏆_�V��G�n�EQ���~�G2	��6�=�[%��O�����U�H�=O��}��SjC>��z���˞x��d~;0w-v�6�.�/��E|�%����¦�^����N`G;18Q ޣ�d�A�'��V��nj/ZTcՙY!�{�u�)�M�saO5F������v�󐳲A!R��=n�$s�z��������&TH��a���
X��4/�SBp�bM����n���BN
��`��p}q�VCK_���������Vk5<�Ά�n{�o�ex�?o�|�z��2���4��݆�\��#Irٹ�4{HL��6��}%�=I���T	� �|�rz�Knc+�|�sswVh@�*c��نY�qƢ�gq�gx���f�Ę>��0����W�\�|K	��1U/�D�4V��֥L!�S:1���"�V`�#A$�*�)_�,+� ��災8�0���Oz������/Zo�a���e�g
��p���r�� ����.a.���ω��25n��w���Oz/��a:j�ם`:*�l��.w~�D����o>�h�r�c����$��>ȁ)��\3��'�Xb,��Ӽ���y��y+*���gg�q�$�y�FYc{�U�[�M�����+ݗ]ӑa��Zj|0���DI�~F����˻�_��y�^A:!B3'��p
���TOzP-�[��
��<L��(��l|��ʩ�	�6�	�'� ]���19�K�B��'���KS���0c[WA��DtO���U�f�,Ľ��)���&e��4��M�ǌ�Nϟ�羆q x�u�[�����F�TҀ��a������J*�4 �j�d_�k�}����x�;�E$�t�{H�>�K�P'�X,���X�5�fQ0�����-ê����
B4_%_��&��aY��wS�D�;ب�'w�!$a���@������ɱ+k�:N�<I� �$Z{��>9g+3�
��yO����q��3f��)7��Q귘�g���I���VA]���@�N66�+�/�2�������S{~*���*�{P	v��Nb7I;_�N�z[S�����J;����j`���RC���T�޼����_� Lg��'���R��faQь9S
�0���<����o�c+�i��	hKj�	w_�6��+Sm:�.sg�&3��e��X�=��D��@s]l�Ӽ��N�r��!������_��<fe�2� 
�����ݜE�(~/���<���W��f$�?UY��ޮ� h��^�ŏ&񸇶Ȕą1�a��_����FlA`M��\t�k�ޒ���pգ��{�;<�-QF sv�N�m8ҽ"�r0@��/S``��W(B1G�5�L9g�����̧��WhG�k90����@�Q�FJ�m!kh�P�Β i��l�Ϣo��B���� Д���=��lz�a�8&f#;<_�^�7��t�&�ri�A�����Zcһ4�����n��5h����w�B1<]*��$�!V9;�׺��,��,���$����N�K|����F���� �w�|2��xO�Z��zd^V�t0���v���3��^� ީ�mGAW#��x�~�����~�h���H׹��_�o#�'���sI8&��=&��D����eF��`��F
`&k<g�}���6V�9��a�lt���[��o��/8��aá>[���t�Z��2_Xx��-q��o����i�eA��z�n�������q��0�\�Azo�lsx�[�� <�������*֑EҒ/�出�	�,��p���k�Bu��Æ�+�(���kȽ R1����"|R�6���j�O�r��Y���.����[�E�9Q����n�����������g��,��Y�S���OlW	~���8�Tw�*�,�9q�$��9�Ƒ�ըP���V�����l�Q��-����p�_�l T���M�C!�FU���uhQ{J���.z6���w;�ة�&�ӿ�my�n��kd�7������\U ���5�خ&軴n�����9�ͨ��$�`}Y�Bw����	9j��\��7}EruM}&zc�W�8��'@O�L"̚!��C�/}Ϲ @da{p��ș{�,�#��@�y�]�3�R	�.�+A��G��PA+F����,��0�G�=Q"�����D���c����*6��e����{�i��
��ZURg��b��DO���d��ù�8�Ӓ�OJG�m���n�ݞ��~c�y�ȸ؍�F��]$["�b��uǗ����Ȫ�V��M-jN���[��e�:3�,M����>��ׁV��o�+b~��^Ϡ��dF��1��u�2z��"�µs�)_/��t�[�qc��du�]ә�����a�ӗ�y�ui����=�oN������[��Z̦�H?M�]9��@��?�	$!=�C.,�C��SQ���<9�Џ�� �t�p�P�Ď�W��\�s��z"��nV��Q	��S��n�`1�Ѧ}[��ϋ�Wv"�[8t��dn����F�q\M�{�L����4g�V��>�<�f��j�����-����r�I��Wc��D���cR��q�*nòY�}Tɬo��=�mϬ
�C�usY|ED��.HǱ)�h4_��w*u�y1��%�!���������ex ��P@N��� 9W��$��D���!�I��p�M�eAh���!~وw*��%nR�p[1���v�B���o�N�^�%w>"�Dѷ��V/�T/b�M�`���}�6��T	�:f5��f�=��b��P_���b��J�K�t���i�h������')/���#_\y�(�50�c%ܧ5 py�8"�<�Ɂ�hH�S����K(7rQ��&�w�����|��1�M従�RL�k���4O� ׇ�yX�rVD3��p+���zU��N:$.0>o�7� N���	/&�E͈�d<]Ev'���`�T�v�]��f{���@�����䀠C| ��"�4���Ɨ�!�Y ����r���W��$�'�c����-iC�$��Hr��;�cvr���<"T�2XY���BD�J�L�4[v�R��Ɛ�r���-oU�M��$�8|��ku�$p���{��s#������gĔ�$�����5YwKN'�wӀB�I�R�h���s�~R#Q��tأ�U��AM��W���Vf�t.�W�\�K�����!.BY#��h3H�\��*^9jW�\>��W��^�/�� �PuA�����A�wa氒����<P��m^� ׬��VO䛍��Lׁ�0*E�
�tNqm%��Z��3p�>	��yn3
�L����nxDW�F��x|y's(��e)̯o7�k(�K
�:L����5|o�=�Q	��N/T��n���K���r3y�Uח,�1����j8e� aE��������p��N����I&T�֚d?���!����e�ķ��'�a��U�MT{:����� ���d���_�M�>�ޟ髆Ŧ� ��z	�r)'Z
M���h4:��Q���«��;��\�\M2���r������D����xK�/�qOqhJ6��4�꯵?�ӿ7�q�&U�K���Im"JH�U�W%�D��2�>����&'nPQĞiog2�.�-��OU�}�o9�u8
����?���W ���,pZ� ��Ȑ��#�u����ZL4��ޜ�e�u�YʬF�hH<1y!�0܄�F 
ד>+��)}��ؗW���U�����褷��%֩n�|�'�=8[���ݞCR��d��e/���К��m��E!������v�d��λ�\�ܛ���u�2&2"A�������b=چ�tZ0��~�&tm��gi��^��3����mQm&2��%�n�f�Q�V��5e�Riit�	�H����υ�FRF��I1N8��Ǣ�$1b��"�7N