XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��FX��i�M8Ŷ=��Sca�3dU���BU�8X�&!�ہ,�ٙe����u<v�����~躧u�qT�Zd�|��2�R����f�m�N8B�#@�@��fǋ����Z�[<l����(>����a��,bѳB��1��"þ5�|��z�y�����9zD.}��Ϙ�W5�?y:N�X�>[?�-�h���ƒ�.=���Wf�9����>���=�8Q�S��_\Q<(ҁ�������o,�}����X<�� ͺe��Z��b;�'�=�B���5rvh:��F,]�{_c�����8IK+�#�C	Q��*�����y_�L|]�LB������	@;�5*AP_��"� U�ϸ�.���ns�ɀ*��J���ձO6�P������u���_���;�S*�	�RV��� ���+6��CuY�t�d��3q��+��Ύ�qT2V�^����:�\�4��^	���|��˗�F=�)�p�ފ͐;\{��Ft��?� �(M��Fb ��'��U}�9$�)Tn'Ǔ��IԚܑ� ���@Y�6��j2�g�}i�A�֖��ZqK򼠔<�%K��d��eQ������`_��Á�G+�����,���ĳ�>&Q ݾa;��n:����zˠ�/�P8�w����!q&����{g��Y�,ܯO��hI������o�&�&XkW$�����ot��5���?�;���綬�H�@�c��`��0T�����sk���XlxVHYEB    95d3    18d0N�H�-��Ř(��6�Ak�%"P�h㷰m�H��~$�i�^�%(m���ur`v�rl�yj����������SFc!��Р����lb��g�Q	HCi�ևl�4��l!al�b3�<���֘0Hޕy�����"�m���$Ԁ�3��J�5sU�f"�ȳ��6�'-�g��Ś�)1�����Ap���;�E�9��p�f��N	qt-���0%MT����4��R�=��l��	s�*��$���\!s��/���7�W5*1y~���2��@[����G�nʹ��I������]�w���aQ���R�s4N�S��,q�7Jc�lx6�!ሣT�o��ֲ���jp�
�1�����<_��c+6�	������+6득�y
�\U��I�i�(?2�
��=F��a���*��fs��pq(Yj��H�P��R�fO0^�>�p���E��@��R{Be�����%4e\�IL���lr*�U��<F"�²�k
���}�w����	q�1�R�2v��N�|�PL��7�v��cu�Z!Et� �
�(��T�g�ͰxH3�e®�<^���	5W	^��Կ͡, ?�� ��,��S��mC����h�k�'���ֻ�;�7r<;�m�V�0�7��j|DȽu��s��C��ǰ��"}a.,(K�����U�Ao��1��$~z�x���e��<�y����O�%�ć~�d��Y��q�� p4����2�8`���g� iS�Q��_���Z����[%��'�.��z�Mp�@�C����y}h�G�m��I6#$� �~�ih	m�OU4'�z���4�� ��3s�Q"�p�g&WC��vw��6#�����Ty����\t���Ga��iU23U�T}�j�e(6~H����6���q$}qǨ�D�e��%��-]�ph��AI �eNƼh���m��?���v��(��؄V&����zr�_6���� �'
�%��*<�'��2�$�Z&�)-��5us��)�H��qȷ��n����oNt<�(3n}kt�ya��T�#H6��
��R��Z�n�yo!:Ž]7�;��a��YE����
z�s6cM�U���rҠ������c�٪<�������\?g\�s�p�(��X�"�C�eY���B�\��6��
��Q*���s��2 h������]Ȣq�]��Cx;�X���Ʒ��g�稜
���ns�v���7���+�7�n���$Z�}7ԄIg?��Q�dS�a�r/.��ui�-�
2�����^�^�����>��Pܳg��9f,5�2A��8�U[?G$A&C�+W���΄��'H���
4iG_ �s����ҩ	���MS���bj��z9��?�z)�b�9b�K7a#tļ��I��.�����m7+�p֟���H�@ՈX��Q3�^�����;���t� ��H���ij
�
Q��3E��/_�G]�Pp��悎%��}!��Ο�������S>l�����g;㡺���?���v���ʄ	2�r��H����2�����ao ��3���F4ǒ��E�Fr��7t���H}���bf��_M �of�VЪI��z1�ߦEX/I����;XʦJ��������=-l�ǜ��o�	K��fO)y?і�d�Sg]fl�����gD���殼߲���B��;]7�P?Z��{MhB��q
c?�B�:������cح$l�Z	���t�Bg�E�D{AQ:V�]�!��6�+q,V�"�^��YQU���x��3A��\R�(�����,�@�v37�ӟ�W��"̨γd�����!q�Md�����
pn�e��nx��N}���I�LǙ-���\��71	��8�f�����`���][�-��4o�{�;~]6���!�~��0�|�ά����f3ե�N�,��'O���ZR~�r��Sʵa=~lP��ɀ����4��{̈́�|�F���I���=q,��u��#d6|'޳Id",+Ԏd?�e\�ŝ�^���B��3$�ZLH-�'�"�tY4�]%��A��į���j^%�e��Q�M1�X��$�s�r�L�N�?�-n��kQ�.Z?�dV"�9(5�;�p*�6�3늉(-�:�)i#g¢��bmPJFA�����3�m�z7�y Z�B�K�Ψ_ٯ�X��3��Os<h�vu_��\�mh���Y�I��
���������>׌�� �`�ϛ��Ԁ�SjXS��BP�"�b��S����Q0�(x�d�b��J��Zpz1h�,���񂨳<��,S0@3/�)ѱ���X�z���+<	wIy�ѓ!GUFo�JAu֗����h:
:%&P�����0�7%�gk����p��?E*K3��R�di<��UŞU�����ެّ�ܳ��5d��d�r���*o�x8V�-a���`W4�]i�F��!@J%�7y�@��2TwK��~ĝ�Q�Hk�h��%l��>�ͭo`R@ 	�=�uS(֕)��6��������㌸��UȦQ
�K��r����1
{B�Ь����7�k���RU��(��\��e�~�a}s��0}q3�$�2#������_C�T	�c�,�	kƇ,�z�j�Z�T�k�������:Ӡ�-M�}��ࣉ�eb�a��N�[�� у�M�T��<��@w�,���g�\�[r~ɫ#���+~���-�&���.&�zq�f�����D�_�L;a �du�h��\��Q	nY6-�iJ����!xP�
ԅ��F,��P���
f��e\�����!3�^�A�7�������K���A���a��;h	Z�a^&e�O�&H!��BGwY�����M�����Ap]�Dw���`:��5���(�ԎK3ܕ{p�m�%���ٔ0 �J �;�ȗ:,�I�\6�fq�g*�@�^x[���2t����VӅ�AJ����1�_>�:�~�OW�o%��*�?��@�=&�s�F���1�'�<�g_�p�HxXC��^𠴡���r�xG��bj�.�ՠ�>��K��Ɉ�����.J�-gN�H�<��n
3��";[�\ç�+)���`�iy���``�iv�C4W�\�*����\�φ��$�#h���ڛe��8/��F����y5��o�	��~mqH�K��5�1�<�4O�Ra�)Q�ܙ�|.�S��5g o����H��| >��<@a.�]ɏ��1��}�ؘ��ze�3���+�,^KcvT�ݕ�
���k��@�����ġ]����#����K��]
_��4+yuK����a���P�P�<$��ғ:�e�bY��$B�>�f��©Q�W�(� �LT �X���
�0�҄ea�1�W���ۡ����Ys}nS���؅�a�U'u�V�2{#�iN����9��q@�%���R�@���lڇޑ��՝��*~�V��q̧�ȭ�{����SI�����4�H_2��~�V�nU��\�H%��B����(&,�K-%�vZ�|7Zb�K�7,�(�ݠ��R�[ʄ&�5��.j��rr�^�L���*	ף�gJ5�q,K�A���ɲ/coq�x����UC�à��A�w��'���c�"~�|0�B��'x��ǔ����7%�
�B�� =�����E��vo��g7At�z�q�\��-�<z��e�V:~��3� �=�!/ȷ !�Ե��c�+p34�@�j�w�I9��E2Q�fW�N����-��B#��c��<_y��i�<MO��ԇJ;v��" #��L��.��q/Z`���brT!�8�&�WAh4�����<�VX&<�O}�R:���Jw��fbjtV�k�6��J���+�U8�ߑ��]o+�Y�a���I����:xZJ���#7�������<�?��.�)��f�/ut�/���F2�����V�*N��7fz�O�J���b��
?F�Gl��q��~��m#6�yL#��yy�[��T���KE��G	�ug\Hߧk�v���;���N�����2�[.S;�R�hFQ����a�yk���F8�VRg����a��H�014�ae]�rbW�� 9ؖ�nv߽ư�t�t���en'�(�SKL�{?C��w���9l����j~��q��8��q���l��;nl.�7$�2��3���0�w,i�߶}3���8t�e��t��6"e|�p�Qe�����cxI��2I�dTƪ�O��� BoWR<s�a7Z�GNĻ@�ٲB[�Qv�����{�$������S0I}[zc�c��c/ƏO��6Y<��H��K4w�����N�j�?����k�@����A�� ����'*q�-Cc�C���(-�$Zd3��V����d0o�������ηje�=K��G���.r�jN:���a��\=0W��$�]�\~��^Q�����pPL'0�<!��F�Cvel��k%�Y��SF��u�C�J�yd�:�(��V�,����`D8`�r"�$!Y���)=x�z+'�^T�n��g/Fw%��K0?�+ɜ/�/d�� ݑ��j��JBjF�),���5�Oa�-�U�;Z�_��h���P�ѯC1Դ<���
p;b,������%�pm���#�F1��P�K���8�f��H��A���f-ۊ��ɋS@F�@�9Η*�����m�$6����K���2��եL"-9���9`O`x�0��Y��&��~�ER�A�����0�3�2��B�{�c����%.L�Ѡp���bӝV��-�ȇ�t���H`�茕��@	�H�t��~KW����]�ecq��|�;�)��2��0;wnO?���l5�
{"Ǡ��N�m5]�SﴦUvSw�E2r��i��U8B��Edĕ0��5+�a���
�(��*?�6<=M& ž(v�����+���|��3��a�֞��&��YW��4����+���Gn6�S���[@7�f�~�Tg�X
i�n��
)",N!0���h.��I������zL�0D7���
3�xb����1�9��l�l{Hм	�%���J!M8�y;Ĝ�~�*MY��n9ڟ������<<k�
�+0��ь���?�5"��QCD\(���A�6�F�&�]ؠ��J�|��7iKx�;�(�3�6UI���L�9��hm�� D�Ox��jB[�d �ف��j�h6�����kׯ]� >����];DE|�VS�??)�-�.$TP'�,?��Om_р�5�i��xܽ���GNX��]����+�؟��e�X�Vd�V�!;��x����90�v4�G�ao��SfbO�Nn�	K=`5��� �v���Gw��x�����ۢ81l�Q?����$�3��K��j��\	�<j��,���4�
jk�q{�-&�eo��oi@����|�E�Б�#�]�)H,������o�'��1/,��i�C"Ä��"�Z�
hmx��7�Z�*ؚn��	=W}ڽ~�+h"n�h��w������Fx�"H���G8+A�B�>�J? ��-umy���V>|^�i�CW�0y�}�^Sv�Z�y���(cّL��!���`R=/��RװMli!�;c���)��s9�4��2���*�+�³5�鄤�	c�h:�%���-�9�i�ׯ�K�����kuo/��_�)'{��tnI��KZd�^Y}T�hB�(1]�����ҙ����4"��^��̱	�wm��?c������}� 7�Je����xVk�����o�#L�_�)�$�V7�0*�0�ɋ=���`s=���f^����D���IG�ST�+i�S��*p.���]�	C�g�g 5��Џ�c�r�_a<8+z�C���g-��٫Z+��'J'��}OBRox���A��Jϼ���(�p�c���ȳ[S�ϺC�MU6�[��_�O��i`ݣ�)###�R@���iȾ��������� ��ws����pKd�{��A��A�|Ѝ��B�#���ӂ�O6Z��m�(���;8�F�7�o�_��)4z�����;�|��Okᩀ��B�3��j���6��eI%�%t�ߟԗ��9K%�!��p0�} �5����t��r�2�0����EJ���Ȥ�"�[G5*�`k:ȟ��9��c���=�p!��fS�L���|'����SNt�й��T������4�֚XRҕ�%[��IyU�"�ɲ F���!=o����O ��H�}��c�N��9o�rE���B.���UkL*(�l�_[g��Rԙ��v{