XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P_x<���+O&t����a'�����ަq�)U��ۻ1j�C�\�(D���'��o�4Q�Ȱ0q�ƾ��ݲ=�ɏF2E�eƣ;3�*��.jz�b+?Y�a�z�b5	��d���Г���'k<���F�p�H�e���8�����I��G��`�Rr�F��<�b��	�)��sS^��\j.w��B�����-�C�~q�$����C����
�׾kZmj���/V2��@>�Տ=�b���-��M���-v��T/�g�� R��wM/j�BA��a�fH�(� Gj	FD�����ӧ����ʐT�!���O�#+����BO�G��6(�1���~B]�z��(�(�.X%�Q�HL��8� Bܤ�qΰ|�ɘfmw �ЎG�Ed�� =s��.��k��(��:�ne-\����擋^�ރ0�N��E��i\3�y��� ��za�6� �_'�ZBO�rM���/
���y%d#a�jO`g�[O���/v.b��F}VR�/�yEĬ�uܒ�"f���j����K|�w~i:N��hLZ�=���jTT���AV�����
~� �t�� ������k���(~��\�i�p�����:gx�lr�=0����iϙ�}����!r�r'��-���Q�Խ��	�*��0b<������^@l�J�R�w!-��)!��?2a���
�#͗��$ �_�������jk�M�Q��	v��,PĘz��$6��i%ŪE������}�I䯥� Q���Pa@O~Jm5s9dXlxVHYEB    b3c6    25b0e-]r�I��J.p{YA؀��
�`KX�@H�Y���r��>�R(�� |-J0�so	������7�d}�!��,˻:�=	:�S�&�_x-(��������f-�h����\�3+�ӭ�|��ը�w�'�JH��p�T�����&� M'�A���苬��p��R����I�G�w_W�i�;Z�ǋ�f�_�w���}��q��Zkf1u����df\�Wj���pW��zq������A��D	����r�7�����, ҳ�p�4U��1ˎ����R���n��X�$'a)S�AuW2��A(�2Cc�C6�R��57�ݠ>D/��
���/F��ˢ�9b�L��߷��qH'4�,����jI�׭�^m)U�?���iQ�\p~�5�ͭ5�ދͬ\X@n>��ڟ��A=OR��D�.B�wj�GHK�r����ر�/0�@z)^S!�f%0&s���\�q����I'��۞�Ǥ����:�g$��F�� �����;w�,E��:��ʭ�o�g���:��ni_Y��O�����!:�0Uɀ�V1Usa5�%����n0�fc���Y��j�+,�i��YB�v[d������did]=��qE�=M���f1��~�K�sL.���9N�ٖ�Vf��@��>6�p��%3^M6mfp�µަ��͠�Z�{�� ����JR������<F�&���Kv�/�����'C7q\	�~lJ9�-<��5%����|e ���F�#�e��i� �lR�8������������ǐ�Z�5j���d��8E�c-��ѶQ�2]�51c��\�aP����{}	46��	tysM�߸l>	l����2~��K
 j��̠%��8+�K.d��)�?))�O�����bq|E0h����Har��f�={�BA��r��|-\9�9�cK�r�0o��u��Q5>�������.�Ec�� ����gJ��E�S��x3P�dl�}AG�m���ϙp<mn��L]�k�Ya���Q?G1�W,nlQ����p�z������y��cf]��� /{#d��H�h��:��V�)��ඳ�z�KO�=�64�e�O�b���uV�E���� ��ʚp{]���fM�(���&-:j����(�^5��^M:��}/�.Ҟ���t�җyX�E�V��X�A�
k/z�uiL��u��Q-���}M�B[�V�ӆ#f\�rB�)H�\������O������a8���z�F3 c��і��s���'����h��d��v_w�4@�XY��$����wV{y�h LB	�JI*d���0�N�3�5�Hy��'����pƤV�O��tm���������@�dS�f�0X��e��V�=�UC����;�&w0"'J"��Z�/�j�`�~n�C�}�{�)�l�rZ����ԥ��K\Wm�8Ʊ�cgJ<JE	sa�a�X��ZE=�k�G�}
B^� i$�/E�ih��~.p%)²��!�
�U8����uY�ɇ���J��H�W�P[1�Kc'�a�Ko��旭#)��[���Jj5%6U��(<o�Z�J���X�Jƪ�f`��5��,��&����W>�6s�T�����kj���bp�wÖ'���b���FHMrRD�m��c�e�~O9"Wep3�'�gW��4�A�5kƗOQ��'@�Ө�{!�q��@��$Z������WC�r�k��B��(��
��V�} -��~.\^�z󓼗m��V4oz���J,hLa��L�\������'f�q\n\�_ {1W4G��*#Z#�y�
r!�:�˃�����N��(�*P6.A��۝��`�� �3E;C���PQ,:�AJHӼ|SP��F
L�B�Y�r�RbF�O�@ ����i��5����3@^̌�ٌ*LV�!���މ�vOl�Nl/�Q$3 쐢i��t:����\�@��3����'|� ���69���Wh�렇[*ɏ�g��Μ���#�ۮ:�+G�̀0��3�ç������O����Tvq~9�3��w��˲X�[�� �.R�b�:0˻���-,��o׈ ��ۭ�t�t!�ڹ_��8]<�Q�I�F�p�8a�6��H.Nc?�k����*����ҭ1�j�]E��Є �f�(�W��+�:�(�&d�KI�:o8l��C�y�P���x˂��_6b���zN�ٓ�H���$T��e�qMV�<K.���>��t�R�^�~mƿ+Uj�� �E��s?��m���Dp����TV���5�E�m��1����鈬+�_�]@J��v��-E<]�P�	P0;��u����.Հ�| �h �Tn���|�O�-4\��[�&��Fz`�-�z���B����0H��r9I��˩f����2�;;3�k�3��.hh�[V��8C�{����Is�I=j�v儓�<�~�Ą�$����.�����U[��s����!����aOxww뫭�-��+�)W\F�U=u�:2i�>Q��6�s�E�����(���	���*�D�J���1��?dd��[�|����բ�*^�F�k�$@����6>�E@a�܀lomC5�����l��+�T�C!B�ʦ�]�"����l����,e�蹷��&�?�b���(�=\��+r�"N����V��6C��� �mp�f������G��w���M&BR|R�%�4}�Ӏ�A�EC�?�8�I/�������Qt�WZJb�6G��f~����U2�L�ZfS����9_m�/��<��{���xi ,�q����Y�1��v�l:KX�ɼ�vʲ��#jw�\�=�dz��LZP1�/C�%�둈XЖjD�� I/'��aP�n`�nN��iL�Ɍ%�Q�[
�|�1����|�W��B�fv�a�E[$�}jE
8�UZ���R���c�gm�tŻ\�ɸ����P*��#@MwU�;�!x��K��7�8���Ts\ҭ��c��dĈ/��}��[Ua<�f�P�Q�L����]`��.�/���#�]�;6+�Đ��f�%���"#rS'8.m=H�P>i-��F	�

K�=�n�eW2�uU�%Ih����h�B��6�#��� 7�����I�d���_����|%�w㍹��x-������>�`��`�7a4;j'�|?�����z��6��5.;O��Pq��&�|F�_��g��'-X���LP�V�����Z�4���c�!\G�� ތ�V���)@j+N� )�����"Y-�����iouJ���y>Ў���-/�����s�2Y�H1��"�>�̍�7}������ƩF���J�(:�T�)�Y��؀��BD]\�|¤X���^�E)�RUk3�)&���׬Ǌ_,��ƎJ˨�	}���+�qz�԰�V<��ZLU��b��t����,�����K_;�3��i�&�5h� m//���K�!�L��=���<R��k`ǐR��,s�}q��e��U!�X`a�b�+>%.���'��c�T��Fc��}I���N$�Ye��~��ڧ�xE�3O?3)�9ң�[�r�t`�H�s���2z:r��rU�Gz|+��7Q�);�~1z&���+% Nȴ|�9�v���*�Da��bL��~E|�ok��T�0fݚ,QI�Y�[�bH�$o�{}e�]xj׎x��������ZaJ��\���g	�`�����?�x��:D$��`GQ�Ґ�3�*2���h�:�r*E]��i�$U�Aw?9�Z���{�� ��8���eQ�qzUƢ+"�<�\oG�am�yt�ҦE�-��|��OIw�^�.�7�Eo��9�/t}+�rHT��mz<��S����H����9B�}���P������X9�wl�lC_�fi��ۡ(!�؀>XӽR��F�%�1�����U�K�� �����A-�ԯ�Kl����%6���(�Vߴ���CdhVxi!��|x�ҶK����>�>-M%�g~�<9����J��#�\�9��6�ބ�x<-F���0ӬA�;�Nӟ�2ÙvVqø�O��O���,��#nA�S�T�P�D7���3�3��1�*���M� �c��P������[�	-���Z@7�P��K�^�!�^������jq2��Q��c��>��SXxf֌����f������k���Z����&�pW�]"Y� �IU�ZP���yT�-�荂6��5:�Z���5|������{�Q-�����ϞR��Q����������um.�m�bu�4��4He��r&�JoF���\��n�păV��__3;@G	��8B`XmX���i<t��7�:�i��eMl�G���n9=�GhkB�WB�N>�]Wz�Ə���M�$��W�l����C.E�߾������6�T[kR�~:e��o}�	��l�w��w!�S��e�b<w��,�+B��l�'W{/Nm�jҦ)���a=o=�>+�<|)m�����M����O��!.d۷�?�����x>�Xb}y���G�A�+�1�6�f(�+��e�,+��g��
S=+8ȍ�s���Q!(���k�
�cJBG�49�@v�rσ�C��
��J��y������Phs��M9��ې���_��ڶ�=?gZ��_�n���y���p�}<��-;,+��\U��Kx�	�TI�̐�n�*�s��� Q2����ON��ͽ-�4�h0\��;��2J|����/z/5Z���4�y��[�qzX�\� ��taMв�����l%R"Y�ԣ�{K%n���j��%"��/S��^���Ĭ�| �A�0��cN�!�����:���R'�<G�^���+��ua'�70/FH����Oj��i�Iy��R#�?~���&���ʦ�O~���,��[�ēa��͵���y�?�2݆��^v��S�m��ב슬�ñ��e�G�W��*�*Zh���ê��dq@o�ӣ�����OWB<������Q�5�u@Ѝ��޶Q/e0vܣ�F����yFf`�p~����+��#�$�&Չ�W�\BH8��jxgg���>r���q-f��G�*��<'a�Xթ[���n�*�'��J}]ଌ�U�7��+�h��#�|�e�P_�?�oJ#�#�I�Sw(�ē��`���<WN�֌�^L"���`�;<~b�n��2�G4������qH	��K����hIV`�B�D��^��J;� ��q����Y��_��2�5��ٓp"� d�Xd����m�	�1��~�
.�@�*8j�a�)T���\نC��./��G�4��q��� kǼx�a.a�fn��w ���9Py��ް{��B�_c��I�Np��i�����zn��0�����e��g�^�����z2.�`��hT���{�h*zH���T�n?G3�~u�����t�F���:����%��N9"�ǅ��C8�<�\AX���+�U�u�����ED}�:!z�w�\;��k#T��x3�us�y��|�`E���6�0ȅ0��Y^G`2�o��k�O��׸Dj�u)
�����[N����)�!x� �����2m¡�Z�����/e?��n�D\jƬ�%�����EV6Q+?'�@%�c�Ҹ�9����,�G����ҽ�@<1NF�R��$ͩ��ncm7`"QWF�x+��PM�:n����f3Ng�0,)������ ֘Qh�oK��w�aQ4�˳�)�E=�����^Ά��gq&�C��F�1���7i��V�3�^�vi����6���LwU-�MiS�e�,���%��XZ?���Bk�MaD�2 ��8X���(���&l���'�T�0S\'MOL'�H��6\��I����ss�k]��ȶ��ഋ���[�WN��e.�<��g�W�Nlo���"��Z��a����QM�.:��HI��N8{�@�Xs[k�1#�|�7�M~�:�T�ה5���Աbtwt��t����&&�u�����Ͼ֠�Y�uU) 3���i׼}�k�d����aHTy$�����~N�`�]�@�%�;���N�&�^ 5�p���TZ�� �]�:�w<j}T�$:KJ ���s���}~Y�SBH��b'T Fq����rIo]8A�0�8=f~��8���0zW;�,:_�L6ypG-�����>	���X��,rƑ����$���������yfYUOF������b";0CJa�AIs23oe%uWY���V ���ɭ�rO�K��������6����/�<qI��C�~��CTU_����}�Ne�z�t؇bT<xL��;H�C����Ap:^T;C��	��^Z~۲�$�l����Q�j1�FOR�T$�/���#�`�\B��G�0�jq��g�u��"0ܭz��ToJ�����Cg��η)���k���0A�5�,w��a�4�2��Sz�}��3���1m~��"H� R?�gZ�ɖӱY�/ 5�w�P���yP�y��<8�W�-���g��d'>)f�|p�l�^Ȃ�	�X�CQ�g�ѳ�,���=�7�R��W�Pl	K�@�/��Ő:��u��5��h��/�H����}[Ӫ#[WL�5�ˠ8��o�/_H��g�U��u��:��x���ٞu�A�j	k=�%D?�8o��1�H�2�otW��*u�k풜+�3ꉮ�t�@��)E�oR�fv&�c���YhCB�5��Nb� KyPv��6F����<�e�~NQ����aR��?00�|��Z2�9K5�sO��ĵ�Ě%��v�O@�p�hs�fNn7�+���Qd����]R؄采�`De��%��A�P��?H#�)=hԹe�<�ʏ���Kk?>��Aj2��ϋ�'�~��2�b}Bl�7�l�9iX?e6sl3��� hi��É���uN� 9�d�D�卑���ꈯ�-򫆉:
�BK���YO��I�\Q�"��C��h��ְ�ȩn_�C:��'���ta�oՐ�H�@�����ˇ�@^UW(�]4�eW��֔SAָmfaaضis\v�T�T�S\��j	SAm�'�є�����n�d�ٺ&���U��8^dz�(ڍ`Q���G��6�����}}g��$�����#-�QD�@�1�.��Ջ0�P�Tu00c�A��d�[K�߁+�I�!�P+3Gi!2�v]�0_�>k
��B�R ��l���>c*&&�mHC�{/��w��Œ�y�0�6g6�|���P�X�/;�7aҌ�L��ܪ*@S���*�e>��/e��8���>��?A@z��>�,�Yf,������,>���%�V�eL�M�:O|Ol�י��0 �А�����\��Z�-@P�6h��
`�5_�� G��c4
�?�uR�i;.VN��;��K�,�F6�������#R��~��Ԙ��Y�]wӯ#�↬����f��&>�\Qa@�K HgH�[iG������V�x��.A���
U�(���[H,-��'Hp'��v�aҠ�R�-ֵR�Wl�� 0u���������=�͵p$V�"vH�X`N,�		�1S����5웟.U���E��=�aܣ��\)�F
^���9��G�ѷ�`4g�Vѿ����#�ԡ��3m�fa�㰁 X�j�>0�4��_�2�y_-�ih>	�2Pέ�zJ�q_�ӌ��i�'kż4d�ON�m�<7ߍ|� ѵ.�@*.Y���&WR����шZ������؟B=�����A�UfǇԦޓ|�/ i���b�!�,�L�(@���s�m���}P)
���CHJ1迫�۟��T�D��Cw��-G��{[1C�I�d�
�±�y�Y�:A&�wd�hv�ۯ?�(Zm�;7P�� 9�O��$��瓽�y{1dt���Ck�	k������L&"��ˬ������H(� �5R锈UsT$ j�Զ���ǶZ���@v�"�˲�n s�L�ڭ�f�`*?'��g�v�m��rr��;�S���x�:87�,Lj(}�����$�[0�v���`,�J9��i��6+ր-��� ��N���������}8��.��g���7҂�X����d1�"X'����b�k���gr��B�󊴈��D�����$�>����ȥ�f�6oV6	9[
1�,�V���V�y�z?��@g�`I=�a69!��ϺͩhP�^�joC��&�/�T����!�B5�T"0~Q</N�m�ǧP$��GA2�]��7��E�q����>ؐ,��J8��E�'G�bS�Pfc��u�D⁇4m�X4��4/3����g*��o)�B^����GX��DF0�P�j�����)�
�����7L� ��n�yM����L6�T�>�lW�C��A�*���c����Eknԯ��o�Xr9�nK�~�F-K����P�.��C����q�����[�L��������w�������L�I����5�A3��7Po�3���>�w�#���hQ |�V��ԡ#�A�^7���M�O�%��^����"��W}ԥ�Tv�l�[τOu�)k��Htj��X�4�բ�ʿ��l��l�v�	��.QCףUr��Փ6*`��p�v�Q7���_"��xc�|����tN�cP��$�f|0OR�Z>��-~Jv�Lu��}���]K� f�s'ǼhU�B����N%	�b(��曯����Gs%�S�gd&�[ �;�^$J��0��Ӫ��!�2l���*���|��2�o���?�����r(�&˜1i`���U��e~���$�b�|(GJVR��}��-�Zѷ'���^�<F���t�CJK"���	
���
C>���'��X�r|*�g{���~�H ^�jg+�&sz�Ө���4&u�я#���;r���Ôn�����K`��9���_�'���M�MkZ���)��#/�8�ّ1ࣈ6e�i��c^�n͗�/�.�Vѕڤ�<w]�$~@E<��s�$S��,�#ĲT�	}��*)�s&��mϏ�d�B`: ����?�v\1�{�4�ev^VGغQ��j��U�r��lh]ٶє��wڇ�Ͷ����%6@|#DK?C�%-q#����=u8	g�H'�q#Jou.�º޹�{]����1�2ݼ~��}�9�g敆�F{�d]K��u��$�+pQ��L��|��>�,)Iǆr����0,��$L�Sf��ц	�SPm��*��1L��F�̳Um�q:Me��/��*���~i��Y��#i�{O�r8��.�˷��ARi���l��jԉ��Jc5Ǉb��%T�\j6�jh>#�Dwo9�:e��э I��6�3[E�J���fǔ��@���x~g<�瞤4�m"�GY� �� T�&��
��<	���iqڿ:h��J:��e�?Y\�55XS�(��u�l�{�=<k�U��5�c��܂P彖v0�4@s�ɝ��.1����^̛��Z�t�`>�{hD�%�8f�@�r�F�S6%#i�//
��(�p2�@�G�"�A+��Xp�