XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ö�ȫ��L��)�?�,b�����3��et�2eNa�m*�ե�E���}!�W�J�cO1uݣ{�L��|����n��7Ş��*G��� �<dxLj,�<��^X_)�".۠������f�W�[��t��pK�ƿY��
"&�b	�S\��!��DVDp�0���(,މ�����P8�}:�ݩ���E-��a3����Ϸ_�	S'{o:gH"�j�|��3��m^eW3��J�U�-����TeT�ZM���^$f&b����܁W����1�^=����<��6�-�:��>��.T�2)1jMm�ol�V���rT׃ƚ��v��G��ۛ����!�-�BT]��`J�����!�i'��n��\ҳ���x�˸�]$D�Lm��7�˾ L��>%d��D`g&���+`��Oy1H����@��r�Q&,jf��:î�no�T\h w����ׄéD[_nva[�:��g���U
�D�&P��^�PTT\��|R4��C|K��%kq	Jt@B5)Ѝp$@�̬eu��|F�",�o�3fp�L�z�p�O��Ei���M��!u�@��O����4���2��|0���M!�pJ�֏����E�4�a���z-�8�ґ\>T1�m�j������F2!��e"ZI�zth�`��r_�.�
6���lp%h>���-A@�Q���o���6WMݻ�Zr�����
�~�R ���YI9��<i�4+�y�������&�����I@�dT)��ء,`&�QXlxVHYEB    b3c6    25b0�0x>�K�l�����\��)������Y��=�ƣ��g\M������,�Lu�������N��T�w� �O�b���ʙ^��.�)b�%߻7�ǯd�^9/L��y�k�[LI�DV��c� �����aT��*�^�����Z�^�{-rk\��e�wa�2�fmw��
� ='j,���n�K�YJF-{$
^�:�դp� ur����x���ybk�?ؾ�Ek�9+։��Z<[����e�<��$zKj"�JL,���͓_������![��%���*ZO����'�أ�}����o6�]����������891�+��eٞ��%�ˀ]��i���!Ӭ����g���;GN��b������Nd�Q��u�Wv�Xc�3��RQ
X��P��ӍT�����Pʊ= ��[�ܛ�fd��bE�]Y�U� /���PX��$5���B���J�4�X�F9�a>]��Ņ�;�i�upr��/��Z߇N�Oy�v;%LVW��|̥f�x[ lg4�ց����B#& 0M�jtm'�U�~�P� GՂ�]���+,0��K��=м�#/�6y�B���6�S�H��v@�����&�&�!.>U|��ڐm��(<#�� qpx�,J1l�6p����Z(~�.�kx��%!8Q@��'������g��Wb�h�e��"�a�[�*[e؋$�ޗ.m�8����9Y�+��y��K���朘��~�xﶰAu�P|�T�T�E����PY{�R4�=u]����p��	i�򲘴y��e�ZёA��[C�����5_�?���3����9�m�&2_)4
����Ik��ﷶ8�#�P�b��Y{���/ğ�Z��um���^r$���t�$��;���"Q��av��}!����~5��M�&xP�N�k_Ⱦ�2�)3�'��u�����j�.y]�[�%T��<��<����7�Ttݑ���5�5����ߌ�a�P-�D���ۅ���V�8.ٛ��ݷ�����9�'�g����
�z��/VI@G*���77,K��.ֻ~�]kU�(�v���E�y1�?��<'��9�3V�e
ZG���zTz�Q���U��������̚Y�i�\AY"�����3q��7eh����lt(�_�����9��۬{��-e�CR@7���.ɋ�u�]p�|nǤ���C�͕�Q����qL��~\�ϫ	Z��+�#+�պ��'q[+�.�g�)����9��u� ��u�:f�}n-��RIiI{�=,4�	/p��:v�T���D�'�ѹ��.8fH)����2�2ځ9����`��M�F�^e4H[�s�� /�#���Ũ[�#��(�v
���Ģe�"�||� ���vhT�����o�!@0��aذ�1H����IG�3���п��df#���w�o�R��k1B�P�Z}ÂI�b�Lec*��=Z�R
���z�=w(@�w7��9C$����<"p��¹g? o]���'�ȧ��3qP`��s����ߕ�M�����	��]`)����k����9��-���s�<)3�~�G�o����{��.�G��ȉV�@��[d� v�%rƚ+߻��r����7$p��h�k[ �����j��x;��Z�Ǆ5�������=6�yl|�����6ژ���+���&�܆*d���**e�qF9��Ɉ�j��d#�	���>Q&�1�ߜ���I����~ΰW��Ԩ�c1�E�R�4��߅mη��<�
/�j���q�љ�
�s�^C�"Ih���M����5X`@�f�$ı�3HD�X� [lE(�v�����]��v�< )~sNN��ޘ�IOm6M}Х�9܍B���M�@ւ)բ�����ѡd�+l�#�Z�Z���{�eH�̞��e�����Yl�K��-,���o�Xa+x�P�lf�Y����)*�r
Dfv�1�B� �hU�E�Do�fa���-(j��X�
)��IR��\uz���FT��b��C�J
WH��:(\j|��]�ߍm#�Q�f�(\�&�3�U����L�ȕ�]�]���}?�%���_%+Ux���:v���^��-��zy��CMx���_fb�N�_���fi�� (��B8d]��U+i�[���17צ(�ǥ<D��0���QO�niO$E
��&hnK �h�n�))ХX���9��x�(b}��&l�By���~�7&w�G&V��hz��$P��,)
�a�^�
-#�=�:=j����Ⱦ�O�����\����L�z�,�_�}7o7B ���*C.8k�j�� ����2Y�^�HJ��08����wfwQ��U�,#��C�Yި� +�my�ܽ	�����CPc<Żyx�#�ڔ *e�C�-U��]�0�tE�v�W�dH�o,�	̂ٛRw��g"t��S��V'z���.��8Kpn����Ugǿ�|Mt�}K.|��Zk�y�p�c�CKH��Ɏ��Ǣ�]��
5?T�76�bY5)�B썈O$Yjz��e������X[�E�!J���^<�!��M�v���K��ƹ�)�Β���|�C���^���G4�3E�{ty��VkܘF���4���7���eG��"	7�Ar5�v�u��	�t�f�(!�~ �������c՜��h����w�Ѐ{�3w��V8����RX�p���bt��{LOq���p�h�&�(����ޥ	�Ts05��̧����0��	�'�� �6��cQly��복�Ee��V��I��WB���D�w?i�jv�W?�ʉQA��L�Gʀ^������(�N�X�
6jʯ�%ٻ^�K ���������B�ym����Y2�ɰ�_�*)���79��P�� �������iu����ҟ]y���1��]w�"�d�������K���"C�,�GI�r-{F	��|�gt�!�Q{�:�xz;	`��ϕ�u��������;S���mE����QJt�h�[ye�䞑3��T�|�b�{�;N������#���ˎ�}��c�	$J����?�7ۍ c![��3�xc;+n]��Ԣ�s��L�U�G��u�޾S�O�b6��������/����Ȳ2���9�S� ) �Qz{��}Tρq~|����t}x�|dF��V�DF��������������0�+�k
>�pP.���i}�������H�t�{ �]~z������1%)o�F����m׮;+�[Ѹil�8�&S}[�o��B1igE��X� JG�H�!�5滗T\f�)_�d�%(�;�;���@νbft92�Fs�x !k-�`^I����a�ZpsMj"�h@w�E��fMXHi}�x(�;S0��k �L�.ٷ8	����>�#�rA_��[�1M|��EX����pG_���;Imx�����YWS�r�-j+ �ӭǄ��vO���}��*�I<�� �t'`�s\�a��w+���]��b|isb�&�P���������X���Z��.�$*��ѳ.��T�p��ɯ����>��9Ә?�Ł6j���:���(��Ӟ���s����v��=���>K.Z���������k��y��&�DR؀̀V-�S�ܕ��[\(4:GP���K.�ʩ5�p�L�
;��ח\�Bȁ��%ߓ������A��
���6+�r����C1�/���o���:sT���zKh�C6�08e������Q
+�	�=����Se�[��rFd�y)	��c�/��V�2`����*8ly�.�>=`�0S� %:�Q���ӿw�)�f��Y��[�j�w�SP�l�)������dI0��V.�P�K�����:8�ZN�İV���	M`Ƿ$�������ҁ�������$���s1Vl�L'��ҟJ�2��B���;�O��#��H�B:�������@���K�4�C�B�r=֒1A�7�P�T�."�]��pH�K����xL��8n�k�����W{�|}�.8��UC|���>�h����Ϥ�,_�&�q��-w�Ȉ<��[��8���6�լR�7VO�_��&��n�MU�B�U��L���QP�E�>�ސ8�K�"%3�%�z� �\8�\��d 	N=Vl���C���vψo�_���+h
�k&.?�?HA���`xK[��Y�	��9���:kM�j�%���_*���-�Jr�L�]�	;��=����~�4K�͋�+�Ač�J��""�A�&�bw�ۿ�S\���b҈�I$6,�fv1R94�h��³i+��H�h8�����)S��B����5��$���kL�f�Twx"��VD�L����L���Ś�D��
  ��Nd�ip�)�S9q��f.U�/��6��(}+���B�_�kJa!�}��	d�r̞������$9c����K"4����0Pj(�B��<�� TZj��k@����뀽���+��ug
���G�	)�ӻ �/�5j~&Gu� �� U�F������>t3�_�oU?�W�O 1Xu�}���&��<��,N���u�m��|ڜ�j�X�K���M�>��}�YmAj��S�n��/$����QgZSe�s�I{ʋ"$�|�S���.��#�}7W8�������.�n�����`}��(θ)(M��fC�)��3���C}�e�g_�9^zΛwo�� ����ַ''����M���Z��K�Z��;��ZŜS?�������3�͎3O�d�Tbo^�CP�E?�C涭b��G����0V��qY����z�����W�׾�b&>�̉��_I�+��v�NX�`�w�SW������N(����B���К
æ�l>=O��u�}�;�)�٬�c$����Wkw|R3r���́�0� <���兜"ۓ7��_�IN�V /\�!�KD0\��4}6%k�[6�.\��������-�B:��s�ʷ���X�KB��n��n�����o���ap�ew�<��E�H����=��"̿�y�8�|2^����Fa,�]��Y�N����T/��|��-T�������&м;�i�'��d��$�kVq��Ŵ�i��P��pR��������nm<BHk�#voF~-.���5(�ZS7�`�r#z����;b���5����]���)�����BA��������`q�R�5M� w0��hw�]�n������5�:�����ܜ����R�J$�!x̴]r$�[ ���Ld������gytu۵��k<�fPz��n)���%�b/./��1�=<qY�3�W|AŊ���ot�dF�Y����!�&e�2}���z�����0�^	?W��7����s1����8��ى�xd�$�b0��d���!��^�w&��ɓ�f�u�w���Z��ݕr�c���}i`
��a�K�����;�V�|��SnJ�u��`�w�n)�&�>1�tR��7������L� ?��0�d���R��~��������U~(8��ݸ�oSht���q1xd�����4�62�{b�#������Ӏp���� ��]�'�0:b�{�d���3G|m߮�t1������ 2�b�q��t�q� ��ޤ�S~?v��n��%��n6訞rܫGŻ��=�^h�^�a��x�~�F�b���B�ڋO�\ m�O�&��9��1x,��1r�uy����M���%�W�E�ᔁ�)�����a~1����y������	�-�o�Tk �H�G�	.Y���e�p���?�2X�Ys]�)*�P��j�.Ů�	ƙ�Vk��lz?h���M.[�ى�n��g�P�Տ��_9=Z)tAʳ���`��'_��̾��d����dU�k<�D,M5WXō�>lY=� ;���e_����b�F�BCjq\]xV[���l�g���A��t�N�"��j�����}zJKa/2	C��O�Ez}�uZf���քo�3�T6��A��u%
�!�-v�6������}ndn=��8�`Qd����GWJ�Os�S�=r�D�^Y��C@�id�%F�چk�vԃ���0���K���궱ٍ�#A1��5�''�1`o��*���;�yM���O�w�/�	`�*B�W�#[,_SD����Ѩ�b���.hEf�k%�;���vӖ�(FO�7{��~e|	�y�7���z0w,��)�Tpp9�_n�Q���w'Tx7���ɹJe�x�+���a�Gc1TA�#��5��H�n��/�9xKh�C�<Xd����+�tD�6p��H�qDP��v�	�k�����|T}+|R|JGWK���@���^�x�)E��l��߾2y�r�R~��=���m�7���k���h������,���^flDZ*��*ʜ�B��й�)�)�6��f�Ja[ִ��f�ɔYʑi��A7�^%5�H8ޓ�[��h+��o*G|n��"T�<��\�ڇ��m'�(�j5������[e=�Ɋ��C�}�S��n��w��]��M�#�޹��?#��"�����7.ٝ�U�q���5tS�����6�?�U{�d� �.���sCloǯu��p|�؁T�c& >�W���:4e8��P�����z�i`�(s���'�9}����ι��z�e�n� )'f�#d܊��P���Ft���gSۂ
lL;(?��0���HxJ�m���z֟y�,�k��迬��v�հ~$Kc���`P`N��ґ5��Oe5������Wf�����Q���<���(ջ�nm�l!0�u����5�f�b��G�;cD�cNk���J�I���]������տQ\�;�*���iC]Q�w��ղ������x���g-YQ�� (u�lr��JA1�r�e�E���C-���p
�&�l����N�?��l�$��+<]؍��!�DF���ޟ�Y��տ�<��E3�z�7�tN���8/�
A�{kK9��"S��p��� P-&���U�������>ŎS�(-5��*��h�c�BJ;f���a%�JW���uF�G�y\OS/CR��L�b�a������bձIhz�}�b�+F�˘��A�����N+nN�NlP�m��Bd���8u��Gå��_��0��č�����Hܗ-���.,/,�Ё)�
����Y��O��]*�xE��V��9���_^g�vn�������1�� 	����e_�ښy.���|b��L<<n��%Ӹc�7����G�����x�#�ŀ�������.��Te��/�� ��<�u�J'��壸�i����CY�j:Bҿ�R�
T�yJ�'+U�B�����(��0���w�e�N����vA������k���|v+C��Ɔ&��R���.ɆW�y�őd'�9`9��*?CQ���zQ����������c�.fAj�_e�4��B>�Է �w��; 6B=�:�+-b}7A��c���
0�j�Pڠ�����~8A�q���G��U�0���5r�߁ߩ�T�&�/4>��<!u�^ԋ�T��3&%�q]����&��wSw����W��_%�l�:���J6���X9�H���G-.ط��'��\s�O �X�璉TJl#V	��*�(���sS�A_@�V��>͖O��ImS�.^]7(u���i?S�쥳P"T���V���YA̓4��J.�<��U��H�ß`odx�r�x�t��a�I1���Y�-��32F�ÏC�57�ƨ�H���h�����C���r�X{�]��^�|���ŏ�i�co�#�ܝ
������0֥��!�H9y��Ɋa�Q$H�'���~_Cd�<�0��9���"����bG����V�!7M��`��g�[�~|}w�p���>�*AItXm[i�.Y��{w��݌A8/�)d�D(S.�_z��L���V+��d��
e��չ�l�v�С>���.��s���VW��|p><0��Dk�p���g>G���d�s$�Sh�`�$�'�T�R��\�Ԏ�(q�d�8�Q�o�@�������,��l}�GYG��%)S
6�4V��i��LG��u�oi\��ɷh��| =!bsk}nI2B"�P�b�kq~�����|G?���	�7������`ұ	ώ���3��	np���C�����aݰ���a+	��p�M�OE�Э|W������^��ӵ,sIFQ�L 1��ixi�_�jŤ�.�Us��ֹ8��	{�Ё�c}�%C��-�,�]b�pv>�璽���3���U��s��n��:iw�< ����:��K%���t)RR��n�OK�����g`�+~o��%SB�H�8���0���B�>{g gH���k"z�n"�`m�>=��G�fA�)~`�*�FP�n�hp�s�s5_'��e��g���
��'\�C"{BD?��g���TH�ef@p�5�8aYШEQ��a
�����g�=�Q٬9�n!~�~�l�P���ok���)��h�;��)�.��y�g<�ļs�ʔ��g=�+��&�>o�]�|��BC�0�4UE��GVꯀ&�d�l"�Â�zk|M�W��+� �POKM0P?��_�9fE��e��n�w�� >(�v'���}ն~��\Rs�4�� ��w���L#��nn�M������{�,@�Ml\�o��iRP��T:]j�XM���l[̀����;��n+=�
y`m����� ��C�Rt��U�[,Q�1�˞��>�9!���Kp��;���0��:*�$�iP����~ ���,XΊ�s9L�:$'����;�?I-w�ŭr���_��#9�K=]���^�T��_�l��u�(1���-)7Ϊ/����1�f5I����Ÿ��K{�����'g�Mh�h�X*�*�a���?u!e�T	R584���fa]j��⫻c���b�`�A��)�/��Iu���أ��s"�jrݭ%��v0tC2��^j@�7Ґ�ڕ��Eq|�<�l)������5x�
(p�Ŗ<f�N�C�?Cv<��N��#��� �����Z_ʮ�e�:�u6"�q�����/�׌elRy�����>����=��_l�|�/VVl8�ĚsR��"��k#oT|���[��m��j�$�u7ݺ�U �s�Z�C#����|����؈.9ݔ��u��T�$�����<H�_|��S"Z����deѴq�KQJe�-�T<��@r���T "�ڎ3E!����k2Y�5�SG�\[5�h3�,gI�V~	L�ya$���M����i�KA�Y��4�����v��Ƨ�9J�q_D���	�6��I'��s����×umZ�<n�� �%� �6�,�̧�����-3�`��=�%Dޒ�e������*|ZP� Ѵ�MV3�0&ƿ�0���u���S2��ײ/]���/Ћ�F3ö����9�9ށMF˧�e?�R�h��@������&I�8�p���]@g[Ӆu�ٺ���E��i�λ����d��#�V|i�,E1�+�_ �%H�O��g�h�_�Bp'
{aξ �3AC���nt��֗t  ��H���SY)���ȱX������J����Z�*