XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2f������v�i�m�f�nY]���L�^^�{�b�O�v�da(�����EX�ja9�����[�mǳ������G��7?�<�*M����ʶ��`�Tf�R�Dx[���D3+�WH�Vn���S'������zG"c^�&�/�DY��B3?.�����JMFCe�����ì2��?�`�-y�����\߲.0�r����'���K�Ŕ�.L;j����<� ������>@���x��`�!Rt�^���r�u�f�����@���xFrM��G�[I3ʡ�:���^}"3�7c$̲�P��O�I�~����@Ն��q$�[�:���`�c���Qҗ�i�;�Y���P<����o���)�߃���J�9�;Ȼ�ݣ+*q7��YW�5P��,8䫚؜���l��%�c6܇V�"(K\\@T�!�\�B��2�k�!���������]���y�o;v�ƺ:.���x;K7�&�lu�4꿱��h��೾ˣhAy&�$HyB�g���U`�>C���P���8u�0��[A]j��"�d����ZU�<�#�sƪޘ/��&��.�4�#W�5ξ �U���}/H��ͦ��s[�+��Į:o�m�]54G�3���b�b���J �8����H���Sߞ3gޑ����z���S5Eø�=-�3Qk�֛���]�YppK�����П�%Z�Q�f�۩ve,l*�ς8�[�a��M��!C�z9"�N4cv���������%�5���.--�A.9^B�1XlxVHYEB    dd8f    2160:�縃���VG��ґI+�0qGur~$�z���@�F,b�<��i��[jH��õ[�fAm�l	� 
�$� �@M8���8��Q��N{\볚�b��) �e%�������J������W�,�"9��,�ho��뱵	���7g�}����WNo-��4��TR�
�q|.V�<���с��O&�3��M�#������+K�Ʊ�?�˕��������
fu';.58�8c �	2�aNE��j�a4��`����R� :nCh��tI�14�3X*{ ��:���bWH~�x��O+�.-�tF���fu��8&�VZ��_��D��	�cB���P���`���6a�q���o�І%Nb�;�fE��NM�4�)�^���̐e���U^0�g8�LG�w&��o)��ru���� Tԩ�k�����N�qGT��K/�ϰ��_����T��{�����+*��2o]n�3���+��p��v
Uh���Pw���,��[����6�����X����Fs�\r�#�y���D��[_]xPT��D�>3bL(��5Ev��E4݊^��w��$�}$
7ɂ]/	w�[����0r�_�@�\M	KV|GI��i��!)��m_o|J���8��= G���6h?�z��[�RvpT���;M�1 ��Єz��c�o�4 ᭩͜��s�3 5�n�����ՉJ�4 Q��a����7"
,�a4=憕�&�j����)$V%�8�sh�s>p�wl�$���l�o�:;����������eױq0��;N�r��F���	�(B�ś6a�]�9%�^�W�l�D�,���/Y��k1�~�+e�i~	���>���x��ފN�<�:Z�m"9%�L�Bi�%��G�00�m����!���NU�8O������Ru(��	mQ<{��G���SI&0�c+������*&�}�3�/��D>�=޺c7���}��ò����m�j`�V����g5�� <�tu�����`�LRތ���G���K���o��L��@��9՚��E��ުm�*���l%��x�FݧF�=j�M��$ؑ��غe.�~��-:�~�k����(��sU�3TǟP��S�M^S�u�'�T�����V[���"��3a���x0�[�t)ii��|t��+�sW��	�"��x6�J�K+�ʸ�yP4�ݝ��};�֗¯���<��,��ۧ��f��x]�F�vM�L,���}sX�	���3�}'zx�6���l`���oy7�(K�OyO�� Px"1*6M�k�]��Z%!��`Z�2H����܆ԋ��=�b3] �)���|��qr��|�S \Q���QmM��$��.:/���V�~�Υ >/�3�9�.���c��UW��T����t�-q�c�j(�5��b}�A�Q��ѣ�h��_U�s�p6��.���C���BZ!�x�����
fB8Zr�E*"��v�e d����K��HtR��[J�]��RBb���8�Qt�'���{$��ˮUH���Q�34�_���v5B� d��C�r4.1JQ�LM-��
~�#�nQ�k~6�@�_����XӍ�
D�a[�;�6\ףz��W�%���=�i3DF!���6� ��Z��C�>;ɵ�ɯ�%����/��)�Y4sF��k���ɲ�m�`���"F}��jw�y��,��!l�[���#��o�s�1�T�>� M����~�/L#XC����EӘ;[�VU�1(Q�Dm ��K�
�iaz���`,N"�Vg�ZN)����쑨�a�l;�R��N|b��Z����ɭo�M/�/��M���y�+ �]���G�Ͽ�h�ټD@�#��o�2ق'�0�|��/#㡅u#��+��'�_���*c�(�g��8����s����A��N������!��mW����.�}�I���	�F�1��K2%p(��Y�c/����o`�B[
��FmQR+�=T�nӕQ�t$��&�gS`��v6�題�W%����.FQ4-��f%ٹ�3��;��(���̍=�-����_�(���������\�X��l�����O�������<,��
ܫ�(��"z'C4MO$\�y6�N
n
�ՏI�u��]L�k�'K��+�1��XK�떤qx�$u�n�$��*ȍ!B�;V����(|4�?ݶ;f���Z�=P����c�}K�C�[|�ń{�̋{bD���˳s�Ѡ�\����<�{����~��0 x�\C_�+V�j-ɤ�~i�quFdІ���W��Z�j}=��	U_v��w����և�Ճ�	DpqR����Ą�q٨]������[��3,S�ի.Gb��|�{)���4SHP��W��W��0�Y���X4���i��!£"��ĶqW1[�t�e/_l��Ǌ^��Hҿyi8����`G�QB��b'l������j��?�yM�\Y�kd�BȞ �P�ܬ[Ro�{�r!��W�W�|���0iye��g����E`k�"8�j�}��A����[=E�OB�Z�f��xY�Ymċ������T�2 ����,G4x����Ԋ\�8x碅 A)���HФWi��s<IY��v�yu�z9���`F�����̶�?o�.M|��c.�wP�Rw�A>z��uR=V�v���/|�N�c��@S���c>!`-=��p+i7l(n����e�'cA�� ǌ���;tu.U^v&i*GI��.r�Xlt��ۅ�J�Ϸ��7	EB��ײ�������rL����5Zg}e�.�8>ɦÓ�O.l v{�o�.�������)'�(������ϑӌ��$.=��1�'�*>��a*D��	���;(� �uRY%9b�o�⸗[<&+|fM�j3oj!�Ez/m��ؚq���3�����p�ܓ��
��͍)N��$v�����v)�t%�m������?@��������_
Ҍ��^>���̇nt���@l�R�+1�AT6��)Z�xפ������4 t�p@I �QS���Q�c�z*u���)�"i������*7����m���$�:�сY�ZT^(�����]`J������A�}}����-

}+Y ��4MȔ �<��+8��lcML�2�R>��o���kE���2b�pA���бK9/,�V3�J#8��]�M͝����8m���nzߐ&~�Z���8}9�t��V�[s�R���FCR��N�c��x����>�-�o�����rP�$1�< ��O]5��:<�G�r�:\)�^{���5��z-a��vp�!p�z+1�e��=��,?H�zi)�e7?-,~F��<	A\�k��O�wO�<v�q8����3S~f�co�ļwD�D/2����2-=gĄ:n�^e����s�?.P�S���u�+��	i�r��nQI8�_i�b$LlwG�s�cΫ� �O���0�|�� ��$�e����nÈ����ts��/x�}�ċ ���9��*��k���)��?�tb0�X>B��,h�P/��#����g�FӾ	�$��aK3�4�;+��?��X���=��SJJ��v���LZi�d���b��ڟ�xX�ͶY)��H�~��� �ꏏV����H��ͳOl�m�r���!Q�I���<'��)v�dt����W�h�L�-&�-hB����]��l���Hu�*�s?��:kٗy'��"��	�f�1v�Wl��{�������5��Gi;LB�����&*�� �/��K�ӷ,B�e�wQ�c�q�c��>%�l�pS�\�DT��]$��`{��,i��N9����X���鈲h���J�qs;iR;A�җ�pX!Cbc+���k�T~�]
nZ(�.�(u�-���<� XC1��ެ�/��]�KR�]��(���/�������O��>��1�h�D�B�K�PfoO��#��wW
�r^��χ��k������%VL(��RO`D/0�hs���s�66��	�5``[
�rʹ�hj"�sx�X�k-Lֽ�P���suZ���zx���*�z�yA��	>��m�ZS�3 �ߎv���M;���+y.!�zZ�	��^g�����Fν���9[�/�`��c��eY(�v���mOk9`F�!���Aַ��7:˪�l��G(u �$�L�����$~%������F1F�����8��*�a�hY�mQ)����9#U�[+�hf�}}P2K�3�e��x�M����j;�Ċ ��v<��JR�
�����q��[lHP��e�����H��ĩe_U�:
���Hpp�\�k)#��[��D�Z$���2�w�E��D}Z6�T�L*WP&i���&���g���+~B/�=���X���]��NŪ�h�v��AS��
I�?�wK�n��Y�3����fh��OΞsݤ����Fv������(��h5>����e!X����7�_o�L�;�/��(����N�e�c:�k\N��Y2S�Vǃ���1j:&�k���[��D�5�����N#��ܗttH`�-k�h�����?gk�H��f�n���H"5��I������ٹyD5@	S�2�X����d���k��nJ���Je�k�ax/�[<N2�gC�낭�O��:	�����lq���<e���G����E��	~����2?\<u]�(k��5����G��ո+�MX��_�m��)J���va�{�u���0��0��f�����G�=�9�Hɞ��/E�'���-W���g���<����#�m�B�$T���*�BgX����!��ܴ�~kg���{uXB1{��$���p~�8�	K���`���RT��R@�H߽�ڂK�J���OX��KJɄ������^U��`zң¹o^�)'�ƕb��ve(U�	̐j(�s�W�����t���YB	�ǹ]���}!3s�{�T
H"��PJ���`�n�XcgLj�_d�y �]Gl�D���J�N���Y�~3����h�UOo��.1����Y"�L��8�=�$c^�R3��/��rk�9�W�g�ňz��g�@ZP>�����R˖�' ƾ��!��g�+�U��7w����r��o�Ȥ�8[I���T�î���%Kw��u��l{N��߳�!u�o*Y�Q��ZZrФz��(?72%�Z��T�y��̯ްd�nw���T�#��ė �m��q%`4�oԟ��˻k8�
���7�{��GB�4��M.�.O&-2�
�2uUO���%�����9��	�d�^���]��Vr1zh��D�����y�m|������9��F��u��&	1P{�1kc�k�����Y�1Dؾ����7(��|��k��/�HK�h�u_s��{)�';�D��͇P%7�v�mۜս�U�z9U�����-���Ie���i9���$�%�:�?��*����U���[�[�9�aW��dft�s�)�p�&љ>-Yn�)m�E���P�\�YG�(�#�~�d?= �ؒt�ޮ���S����.=ܢz�4/V���:���;<����:��zv��38t���\W�*(Q|�y?h�gdǏSrQK�%gp!{¢gv	xs�0�D]L��s=�)91�XO�÷� sՓHA75F�88�ڞSN2���I���/o�c���<�d���L��+�fh݈�u���z�/_�C�
R����Bd25闗�f�,>�LeR�b�h�)���bL��8)
��K��2��*�U��ƍ��L@Y�^�oY�aM���`��/�jѨ�����],c���^��ٕ��-�!p�g�[�d�_���eb_
a�~k��[���J��l7�{��ϥ@�m)h� ��>T�v�D�2K�fçxL`��{2ޑ�N�K��O{��u;>x[ѵe��G��	A�Y�J��cI�S��K�-�\�m�9$-=γ�"3Gt����u�Ւ[4S˸Kuy/W����_Y�u!��f����"����}\/G��|� �J����(i# �W��*���*J~ߺ�Vu5������\�*�fP�����9�_ͱ� a�Z�ӐF²ȌeD��n��/�>��z �e�4�{��*և�&ȲFWNF���0Ʌ�\&�ʃK0������b�(2崔���H�l:�XN"
�� �o����x�#50:~ĵ����g���5"w�i{U.%k����|�5��>���;�a�;/�.p>�)B�(����/u����#�r��&y�XN�_YҲ�����D��I�i1|% h��|�xo�D(��v���{���
��V�1�����2a$��Y*�����!�Z�(?�����X��:"��Ǳ �W��xGs��]O�|�G�;*�8��pm�葊o����y�;�>T��h����M͑C��kЀ_�S\X9��9��d$��'��~{��ށ��k�o���0��jv�W�6��[L��Q~���X����|�␒@粷�g�u�3óqYq��gs�bV��ej����a��v��X�J0{(��s��<�gN�;�����g.���G��&�K�(��S.���_��r�2[Uow����p)9���)_7q��P��I�ـr>D�����C�J-�T?�+�n,8���y��/[)� ��]F�tl��"��n��M�@��UɃ�J���y�J�4{v)�Ց�̛=	����K��+�cDAi��|�r�������?�&ӌJ�Q�k��"��y5�-F�W]��o�%ΞWBє
Q*՛��Y��Ǿ �5��fX�����Lލ�R���Ҟ4�����
�xiq�ŏELE �I ���N�x�qs.��LH��4t@M������X�� ��"5=�7΂~��7��*d�L�^}�Nv��,����ŏ���dw����5���o$g�H]�xܻam0?"�.f�đ��U!*(w��6t�i ��������b[j�����;���X\�!w]z�З#d}�ի����+���TK!f��F��5nv��)��q읝K�9�>�8p��J��}�( ��/d�H�v�eg?��	ip�6'�  F��!w"DRd��n�s,u���/or#=��)n�Q�JǠw��"�߆����V骖�"c\��T�x�Z)������Q��Py��U�K�˃K2T�Sp�l����,Y�7��`�	��i/R�UO�?����R�(��(�D<�I�6��^3w�
��hٞ��,?P��q��wGJR 0�'Ƨ)���gk�Y}/^�x�%��3��+��<�m�<Yf#�^c����D );��h��v�-O$��yY�L�2��9+�ac��_�G�H,��J`�ցMl���5�;=�:�W�z=`��V���~�ΓN�*��GR���RMCԒ&9���⠌v�\�<��b�*|�5��\�7���3G�"i��(8�Ђ���Y����'�[�]�fĐ�򺗣��!-O%=������2�
NW;<2�%.�ʂɐ7�M���u7N�9��uu_�*DB����ƚ&C�NN�<0��8{��43��F?�꟱*V�͠������sf��)��J�>��@'Z��.��`\�J%�p�5���-��I4�t����d�l��ҵ7�D��8��KQ�,S�B:Zf���p?�L)'<|d�����0���8�EZ����;�3��זˠͲRp���1ʕ;������D)��✺'�s8�'�:
�M�~���R��1	�:hZ�Ծ�㟞��$�|0�t��o/�:'jY��
�8��l�û���ᱳ�,�ZK���)cV��ge��_P OK�kc�M8�������.��u#��JM6��	��:ǳ�C�HeI؎��z�m$��?��E^;��������	��녬��VMY`<��PT���e��e�ȳ�&�v�R,�� U��M]�^�؎��c����Ж�b�_2��;�lZ�$+/���l}s����v�AQ�w��c��`�����E2v!�؛�uE6�Cv(pP�I�������mm�'Ɖ���O?�q1n�z\s��sݠ��w�O�����}�Ձ����|Xd([��H@|}����<I�}�Bd���ilƠ^3�c#�=�����
�zT�Vs����`�G�bz���?]�r��a����%�������{zϼ�Z�FB��͍1ZC@�z*Td���M�еro~7��,��d�l�EQ�f3,��_'��l��.T/�dP� LH5��DR�@� }���Ld���?���;��|���x1�'k�x�ω����M�vа����
�i'����2�ǔvS��� �ve�[_�B�Y��h���5�+�<�q����0ʸ����@:�+��ʶ(�3Up��(��;��v�1�7,Iٚ4�I9L�8���������HLLOJ�?D�/�{J��@��: