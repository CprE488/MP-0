XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w�N�C�#���V����&a�D���s�a��(���{������426��[;�i���`ik��]+ؗ|+�@� -A�s�i���!c�?�+�l��kH�~����A"�y�l�8(��B�{����fR�E��)�n�- �R�n�N��j����=�k籏�h)�Ye�_��U�tu�x�^| EƲ��{;���K�E��ƅ�Q�;�^>V�����
;���'��Lg,qbЂ�8�߾g	eM����� ��0j��}�RRP�16���R;��J.�k4�%���Y�V������a_����.�{Wr1e���^���v��T�Ƴ ��.D�.�Z��a�����ʐ����x��9����_�d@1Q]օ��3����vЀ���i�}^�uɵER�%�c��l^[��4�^�����Z� �t����{�(�,�y�/s�=�����4��x�o�����F���c��T�5���H�J5F�䖻'%��C?a<�7@��/�"`�I��@n�.$�jٱD	���/6��z�;\�����u!�VH�t*�U0]�۽�ކc�yt�p��<!|�B��\{���zt§J-��r�SV�p�T�2�ْ�0��i��A��N��2�5FRrž��i+��5Ϭ�L�;e�����Qԕ
M��;��� �8�x�y9��MqhIL;�����z�+�ğT�w[v'�c�EW�{e�7�;ba��G����5+�$J�F�Jpd�LӶ�gp%����`u��~���AGd��G�XlxVHYEB    42ae    1110K-��?�	#cx ��_qq,���~�!��\$ O���H��j�(8�VS�+�� ���H
�d%��p�~0���.������[�{���9���E�{e�>�r��=){{V.'���p���� ���A�q�d��Qe�Z�4�f��^>#U �ZK�˔��1��,ȶx����s�����P�.�=���2t��=^y�M�������2?����*;�a�����H���W�a4שy��|�3b��qM��J��d�K�V�e��⒪�ș�И��=�g��p��]1��d�0_ `!BX�	u�%6-r�q�N��D�^��f�j�=G�~W_)��8\!As�3�̨�u���td�d��ϐ��W�ȟ��w�.���V��N�_|3�bp���^;��-��˯qN�Z��O�/ܑ��g�l7d??s�����k?�e�4�Z�Tω��Ig��zy'r>1���M��v�@_E[+X,�1P�����\�u &q�F��/ft�nxC��_:с+:�)�����i��AGc�L���yEln�1K����a늤�Tm^W�v@��uʼ7�� �E������asRK}!��k[�� ���s�1���C��&N&l���C�X�r�*���}g��T�RPt��/��5����P��k�6���U�P�2$���Q��ԁ� ����cOǗ#v�=OΫ��2�#�G��v�CnKٖ~c��Xe�q����N���_e �6>G�ΝԒ>�K�M��Xu���X�':;��7��������~���� �����K��4�Ga������L�	2�0�r���Z<���<������-�����5=D���`����`�4Rj8i^ ��z,��U2�6�e���զ��7s`�0�������g��fT�7z��#��� ��&�<��\�Q��!��,O�띦/���!dF)[l��N
siE�d"1�����cJ��}�X&��~ҵ2z�z���B����fpFd��c��q�t^F��U<���5]L��|Dm�"����}3!g�߇� ����۪�T)�u�S���)�b�Wm���FX�:w�*Ω�������fo����sw�*���?����4���D����Dm��aE&� ��Q�|D/��m���l��Y�*z^k�}Y��ǊTOu������JT�9uB6�[1���/��x�)�U)�z��9$^�ñ �oೊ��f��Yw��?�Gn�rk7b�����Ҩw�|6ȃKn���!:�������&W�E���3������X����!���<yS2h���bSA:�֨(~��);��p2� &��5R���C�9U-�D�c|��H��~�����4�'�T6���������'�<�7���C%�;$)'��ڨ`�H)���O���Ҵĕ�&������*�bv���t�O{�CKa��l��
"��MZ,���W �j����*D&G�t���J_�1[u���IJn��MqD�Ê��+�� {���Lj&������: I���S�^�fΈ��O�`#Q�}�a�B�ᤪ���WN��==!���^d~���F������������@T�hmn+�+.� eFs z̅B���G����*]0�.s�6U�FԊtcZR`8η��[q����vw�������z�v�����3��Sh���hC��Ȝ�C�N���sþ��\��	�Ze�tӮ�E�"mL���`�)MF�1����Ѽ�Jj*�@�D��jP�Rӗ�K?�∍U���L὿�����![�鏲C�jk��Ƹs�OrV��<��G��]L���LY�7CN��0hИ�R��1�X���rT�@��ל1������~�z=t�YG��_�x�Pk3x�����Ԣ"�o��Kِ2����4�:�r����s*R0(�_�i�&e1P��N�g�لv(n.=�s̅cFWek�O}ɂ<MG������?:y,����B����qF�����t���a���v;�y%ƨ5��MPNgȘGc�}egnd�K2Z����Z�
<@���b�B��g�SⓌ��d�yK� e�RW�0�y�M��l� ��� ����&\��6A�p�3:S����s���zf� !��&.�L�U��2���,I���L��tq����5r.����J=)^͎]bnk|�5��p�	����WG�+�������L�;�ZU�S��=������S��%�ژ/���lQ =�����Ŗٸ�)+`|nl�������(	4R��%0���7DF�F[�dME@b�����g�/���2fg !bpI(���@˯���B��4����T�(�p5���R:d9�e�ٙhn��v��ڜ�6Hs��ȣ��7 0��j�F��;��_�4�����]S��d�H�s�s���,��nN3ֿ���;������s
�4Õ.�:`�Ce��5R��}��Z�TK/va,r'�[�;�^j����2{.�)�[�e�U���V��М?]}�%c$?�mh�hX��W�ǔ����xp��ǈf@`�u!>�S���Ի�m`���/�9aה�f�(ױX����h�g�?H�5�hx�������e�[�Z:,\�x5��L�L��R�9���)n����*��|�s96��R��"Ϛ�V|�w����h�	�Q1�L�=iK�Uc��VdzaI<Ȱ���'��(M�4>�����oE�5.�S���U���L������X֦Zj��� X��\T�A���GS����8Ӟ�]@�N�D�$�����0���>0[�:3/���d`v�ӏ��P�-��0Ɠ�`�n؈�G>׽
6C�}�]��\gʹ)�[�W��Ԁ�u,/���D��]0X`HI?b�S�|�� :�H�x�KG�k�J�
����n,!�0���z�6�;���D���:��H3�99 2���H2;�UO>ge�G�Ä2��B�ǀ����q��F�J���{��3Y`'����0��e�x$@s�|?T���5����(Z����U�J%zE������V�.�(e����ռ>��w�C��}�����c(������tkqNp.���82�����Z_ç�Ѓ����
IDf��q>���&��Fb�V)v���Wc�����9X~@䂻sF	\�3=�}w�q0>=ʑ��m~ٞ[�l��ojT�boM�g��$ۥE+���I*�ff=�yrf��������Q�ZNסJP��j��o�Z���({c&�=�s��{ dc�{]�Z"�["J�&�pcB��� �nf?���D<��tqC�=�UR��F�������������mu�Նv�����[��U�ⷄ�D�ǎR�Y������e�b���p�e,��p �]�Ut1�j���o��@慡�Oo[�+L=�����Z
��]�񴋷�i�R;�H���w����3I���/��S�Sfl�n�غ�]3`z�y��={�:����ME�wrB�礽��=���O����u�ކFY����Ks�.�-�g{��H0A�� �ث*S�{���m����0�un�:���djYj449_f�w�@;�fA���O��5�b���K�Le:�(ϲ��3k�	
�����/�L �����C�<���<��?D��ƄN���_?����+L��W~JX����G	e�I�PxeN*y���fw}
��d�s��Ni���O����;6@��D{fj�9�
BB����pL����\��G��� �r�������3���m�Ά	1���^8�h4�^M8�%jƮ���=]�(��w}R0�czr�X��U�8)���E�QL�������ց>3�5���o��2[�XF���:9z{����������L�$6|'��"U��8�:�j���Y�GP$���Јo�W�G]�2^������s�u�$�m0�/K0A�����z�X�`6��3[-���'�O�P�!c��xp{h����/n��A�{Nmj�E©�8V_ߍҁp�c��ЄU �.��2�B_�RJG�ڱ�����̪e	�ryW�Q�w���Z�[���"��)�
�脷����,�7�g9�9�|f���{�?��tb�1gv]{��T6C5�Q����g��&a�*��K�W|�sDkI��¦ �[��7�Ojs�o{���~�ݡ�r����aP�	XVEy1<�FgLP���v�m_�2K�L�ـ?Ã(sPG��