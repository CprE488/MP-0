XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���=1G擈W��~�K��1qa��cu�-1RY�Yb����&C�[����/�E�*��N��uߪHVW��JQ9�
?�C��(ʤ�y����v�%������̧�,�Yrio�g���*ZH�ld(%oGG�1[�F����3,����������һ�A#df�j�g^����1�X���&��ve�_�4�����(�6���+X��Z8E0��N��}u1!�g(�������HD��7�2-�a*Lr����y��r�eS죦>Hsܩ-���ٍQ�%�q��.��퉳!��Z��0Ǘ+\�=�$ӥ�cv
�r0&[�4�.�wM��古�VG�f'{L+��oMS�����W3��忯���P)�:g�i��`�0ْ��:
U�D�k�f:}95b�}Y�qG�ж!%DD
k��b�N�4�1[��6�~n��k.������6�ߎ�<�
�p�U�
�h�~�ڿ-�\��/�K��&H������`5�U��M�|c���]w�=���H�uàBR�^�t���?��sa���b[P�
��9]��v�`�˃ty��\���^� �}�%_�ԕ[':�ٞja�Bc��&C`�@u/ J͵S���S���K�vжXj����R.$lV>ۈL*�Pn�^"�0�ǭ��o&}��/��	+'*���;~�-4֛���(����$���x�~>��V��n��P�T�O^��z'i����B�y9HJ���O�XlxVHYEB    b3c6    25b0�/��F_��`���I����a��¦�aU��]@���+�;6K�K۞�9Bd�B�\������C��)ov�)E����f���ѥ7�ĳ�G�i2E0���3��4c��v�yfwe�p9��B�/}��BT*�WK�x"����), _��n�	 f�k�KѼ�1r�{�V�E�Ioͷ$�c�#K���Ä-������``b�� �s����,�kt���q(�P���O�l9��(�������T�c�\��!� i�@��d|�7���k�g7���w�zP�Iz�.
W�d�N���=z���֭OPr��k>�x	��/c��;�<���W� ��8R6@{���B��	/���T}6˄��7�q�K�< )/y��m/�_v�확Ӧ1����|�Y��l��c�kE�p�xlv���Ld=�`O���� g��黑Uŕ�h=Ò�Q��UT�&%۪��Np�ٕ}A�s���(���C�c��rmM8腉P�P\��S�q��<�r���V��(����,~h�&���5K2� E��>>z�4D�O�l�AT��7��Q�?��ׇ8���r�v��ji&�W���l~�Kd�7��Xt���4V#�����L�gZZ��54������cu	JN��{�*>�n-6��.�4:-�`O4|M�����j��a>���i�`Cn4�~�f��]����D��kqm�[_�v�/������_���b����U 쨻��R�b����-H��G%`�eN���#����'O��l��ߧ�4L�C�i^����)��۽w�PLſ��R]~���>=���x64��1~�^uwb,�t�Ur�	p���=�/�z7e۶<0�͎:����P��: ua�#��#��'��˗�R
�(?���(-�~ꭣ�A3��s1ű�{kt\s9s���[7����g W���s�%H�Wg+X���騜+�~����ͦ���'0=ڶ.  I�oڀ�ݽ�.��(Ţ4J�����?���}VIT�s�0�ߗDG%}����E��M�sn�5���Ŏ���� XK�y nהv4Z��n�ʈ�I͇�,	��7ռ��GaYS3�avk�&��/��Dō�F#�ru�r�%�� �n0#$�02éE=u����/<�{u�Ո))��W�s�C}-��*�+���)!R�!j`��.�A�~V99NC��R ./�u#�m�JaW}�W��	'�n,~������,�O�<6O\�8EFz4�Hx�(�rĶ��|Ǜ�Y�cC�<�SA�;v��T�]�5�be,��ɠ�G$��ޙt�����=���e��˘>�4�����s�v(ع.��C���s�?�#ù{�
Pd��#\K����%�6���)����ù�S����7&b��J}Ⱦ@N��p|�!�׆fZ���S���buS�^��B��L��׵��#>�7�����o����JyO9���j�-�kc��?W��W���	�گdjx�#���TS�m���P�����ӳ��}L�C������8A=��Y��E�=�?j��Z�MEsL��z��X�J�z���U�8��E�b��)���TU'��-)���m�!��J���`�{��9ݢSM�}#_g��BI8�_$��ूƮ�)�R`�t\��A�X%�@����n��L$��_�0C�!	O��۸�q��kDn��H��۬�,����
@�3z����柔�у��H��k������F�p�Jr� TD�c�@�t�j�����bk���L ���#�&�\%�2�7���!��0�n��%Er br�)7k��n��I���6���?��J�Ô�1�h�cJ�ە#.�f}�ɬ��������x�݄���ѵCܑ7�.xSZusM1��O)S4�~�iibf��+��M�ڋ�fV4�R�q �GH\T�W5�����j�E�I�Pe�^l;(�{�d!��}��)�"n}���A#L�}#yN�q����G������0�����=����g~������e6~����?��o�Aՠ�AW:�	D�����b�<���u�p�T���"�ɫ��`:��ԡ\�1:<�j(������?)4�T��%���2��\۝���pӫ�A�3�C�F�qQ�y�E��׳�>:�z����$���i�N��b�x[B
�-�� ���,`a��g��	�A�l����o�_J�~��Sh�ʼp��ֲ�v�9'��%9$�Kr�
��u��?Ѣ�LT'jO�d�y"fUG��f8��}
ݎn��F��G�*#3c{��Ia.�f�����p��������FƮ�Vډ0�dZ')&��yV:�����a���6^T�o!<,V�[j��y�H�9�n�4�G���6��d�N6�Ԁ���]�d��TH.}�aڑ�Z�����=���l� � ��r��E���v�{��
~�~�2X�q���RJ$\�����7�_�|#�3��,��_ʖ����O��j
0&-��m&���r���);��� �53S��d;T�ޒ�;Ǣz�LD"d�D��������:66�y�]6o�rP/�X|�j�r�ʍ�ؖ4\�� ��駺0s2�RS�ɿ�3�����9�$ל� �>x#A�8~�w+a5���2Pez��T㬿Z�|�U�_��T�ॻ�Tń�RI�^��j>
���XNmo�t]�[3j��ˡgV�O%,�D����
�=�������C7��¼U�:��n����Y�C�Ђ1�(k`�!pG�f3Mj��z;1�'�i�6�4���5�Kc�:J�0������-���Hk�h�u���{��t-�Z�s�-A��C�WY��-���Om�?.��q�|���9U�n��U�
���P�D�P)z�S��	^t3p�(��ԿF�ר������nsqޅTMq��I]1؆��c-�|U@���M�9	бvu=�7�7�P3?��勈���t@�'��0�i��LZ"'��r���U�����|���<@�䐙:�W���|��RYl9��	��b���g�����3�,��S����¸q��hHsI�G��n���4�K
;������ؓ�r����	)�(�i+S��Pw��a� �k�
�1��!]���W���Pr��y���MG���PUz�c�Z~��C��Fp�+|�yD�+;ߛ�)����n�%D��g�ȶ���*��xn4�2 ��r��^��q���f��� a�+�\m����.�lta�tt�Z��X	c=E7��9	A���j��v0ֺ�F����a���>�T�#=�S�<ABǦ��@�ޟ�[����M��ϫB�c�5p�ʵ��r��a���	�DT�����*|�e�����j[�� �d�
c#7�8r�b����%!y�y�#�Qe�D�����.��лn����!����JR����ϲ�o�=�:X�/����EDd:��Ϟ�}Cs�r��wr��m�i��(��Szf��
���k����kҍn�Y�@Օ���j[wA\�������5�$���"��<���RA�OL�ڝ{t%f�M�{�aPKI񕠘 �dF�4{9�j���]������$�g8�xI��]�	��|�*u�&��9Ub~�8�'�����?f���\���У{u�~�͍����]	�:�}����e�Ѐyb��9�|�L<���p�)-:S�;H��d��`���q�Zu.r�!�g{�+�>�^�g��֗{�O�h������,v�S�u��l�C�傗��i��9	-sX�34��X�9�	kN2���Xt�%#X`�R����FJ������J5n��I=��t��G�KD����L�&:/p�� �4a�j�5@'�-�n�7�{����U�u�$�,K�;�ĦPX�Vb��#7�_��T�QN�C���_d��T����l�>��u��B�E�i���u@h� ����zC]- �rJ]�Ts�f��J��J'��x��x�W��ߖ �J<Ç»u�r���s��k�&�Li���B�w9�VH~�:��{�u�8K��0}u��kJ�Z��s����E�ɟ\N��LUn��vM�E{I&�,t��B8�)�ߏ�X����2!	A���is�n|_*t����z�s�R�o�(|�|�� ���Jc]ΧN�y����x5���0�7y�a�׀5�y@�l��P���%�:E�"�ca�E�7y�g��	v>�Q��C%�i�L)���6��bE��	�#��)ДS��A�Е�Ec�{ۭOc�J)�;#���%����'��[�a�4��a�da#	Y3M�s��g܄��ZH���)C8�="to3Y�WY����2�]�"���Q+��+?�#�����Kov��"$���oR���_1�w�� i���E�r��h'�)匳.Df'�z:��J^���m���<�M)��a�PzJq�t�O���������P|,}��wFL��\ڂ��o�B��fn�l�w��
����X/=�懖��� k�gcR�����k��5���,��q54O��G�k�CWhT�vRR"�dF�>��ǎ�A�̒O\D�|��ᮿ�a������EA�K��u�n��${h��G�Q���]�Ѳ�G��Y��a��bd�e�^<x,E�ϢD��ҕi���ALHOl
�ǵ➾�(Zo�K�#��y�C��"`R��Ig($ �	���Jmȳ(fg�=awP�s�R.�R��7�Tn�Q���:�{�ǭiY���ܧ{��$�$�T)kb�z	�i�T�*�|O�c��ʚa$��.{���p�Q���U����#AS�Z�튐�h�1wa�1���6i0���2������cJB�D���pַ,��*+K;���(]����nd�3����x��QC7^[g��o�z{�Å� ���`����T+���V� �y�(��~�`��3k��͊����Ϫh��C�K�ߊ�,��c��[:F�P:�Qt�z�\��t�}&i��A�H��c~J�ŧ�M���l��YB�>̌��T���b�V�;�����Q�$�H�N�F�8�����`i
��E���rŁ�y��Z-��^"l�P�u�vmA�����+�W���MS��^0�H�Ӎ^0~ґ��� ���m����<�����F�Y�=��&�v+o���g��إ�KV�Z�6<�[��>��M^�{�w å�ĥ���7Z�O��w5	k�
�а��5w. o�銊���E�����b�S?~$��F���{�:Y'�u)��	+.���Cg�)Y�?��.bU��K��]oɅ��\ $8r_�b`j���m�1����*��}ā���T��2;A���������--%����m��9��T5�S�Ó��+�N��V�È�Zp>�=Nл��槍�*����#J%���q��c�%��͌�&��N�CI �g��y&/�����n���`x�60�.�-�61�y}�p�0�u~��Փ�E���g����t�`!)�omUAde֓G�FP0�hmց@��^J�iIy���`4 F}kP#�VU�]�C���&���R��{��q���;������N��Oj��޺0�P��HY�w��!'W>K�X<��!>�!�f}�������kCE����"7M5 Y��Wu�h,[Xc~w��b�W9��b!J��S��=�O�����ﶒ�J^���pZD�:dёւG�,'a�R9��HA�4����%��U�z��C�����%�L��V�.%x�l�V���M=��z��l�N=6ˁό����;�t�RGS��m�g}�I00haA�k����r=&W����|1(E,#Zq3#a4�0]��1<z�hц��qU��.��r�S��	��q� a*�ښ&�U+\��!��1���PV[g��:S�<����_���Q�O��*�Pg�n�����>ÑW���<�'j���5��j�U8	��.�r��^G��u�
�6<FF��?�7V�F���{P����37h��*M�������eHs,����oe������}�C����`�L8�/_y��2�/W��7�T�}��k}($?rp&���v ���A��DL��"�W�d�iӁ���S��;v��6s�1��HF��|��f��r��u���x�L���fH�'�.ρD�3�i��>	�P��*�P�By�?pɪ���
Tw���]���
�_Pr^x�p4uavj�)M�p$p�i<c\�6�"9U���A���䮶�g���6��.��jᖕ���:Ĩj�P�x���^��Gj@��H�0N�� XX}ɝ-7��>�X5���j�c�y5��l�ބ�<��{�ڤ���>�5 '�P/Ûjf�i)��)���v�n)#�"����$M6]C�_Xrh	�����Y@W��E�0/�u��n�xg���'��<b���])�#�:؋���E�&ߙ�*�ok]˿�k�����<�`����]�'��(��0�^T~�i�D��ޝ�u�:K:$��c�����D�|ؽu����u|T��%r��uoR�hCYi�l�S�ʤ�u?l��[�C�sz�l(�����_�<���Ɨ�Lb�t�6���=�����_4:�A]j1�\��!h�W=�1�t���8�ʓ	8�������"��{?$#��c1��6�ɖ�S�����vk�P �b�?vT�bJ�)U���?t��r���u����j/���%8�O�F��Ow�en�Դ����	��YY��Zu�KU[ߗ�G�	��~��2p1�y;�h2.?7��瀓 I�/�>M�e{2����L��������W�94���l[�ѿ�ҿ���F{_�6�6Q]��+�_?��*x<�=&B�_U�"P��6m]��#|��mJ���'
� l�h�T2�*x�ʕ���Ll�L����dޅ8���m#C�i
��-�-��od}�X�/�թ�s�az�jǒFr`m���@�.�=�\m�yYM4䢥=y��X���xH��H6X�'qG����(1��!K<�6E�'�b���T�9��.z#=����%�T�߱�yq{�?i�'J�}Nxœ:Tk��ov珨�=����Ξ�B�Y���-�GSI�}��f��aV 2����4�}������6�P�����"��,��+:ތ�Ց�*a��V��/�ʓ2�c��}����[õ2�=�Х��=>�\�ֈ҈R��V;�xL�ӳ�p��%?�����
�I	w3?���G�����=��g�����k�o�&ڐ�iK�fDklv;H�FU �.ƶ�y��J�H�"]P1	��cW ���K�h����I��G�IU!R���kw�U�^9��2� aj����R�RE�Η2H4l�'u���w=�r"���|�Y�#�X�ab)V�6���J���Ť/ � �iI�AU�����NdX�/L>��� �߫A��$�w#U-ۀ� ��G��M�笭-���yi���]s���z�{ �#��u���:ӿ^w.&V��R�������g?f�8�7G�b��ڮR7hX��)#�
`���^��Y�Tao(H���3ܽ'3�U��W��$��7���H6V\*]�LW̰C�'zl�j���2�i�C�ts5g���=�s�É�4���ZD��/]�����jA���}l0�H+[U�4Ϥ�[��g�g�Ƣ4���:��_�h�X�d4\���˻�~J:�YW��o%[�<���,���U��:�k!�~u� ��X��t����������l�����d<�>F��6i b��5�K�0xH�L��]]%�|J<�XC���rBXB��0a�Fz�c7GO�l+t�Ѷ9�N�������$���·���=;�g�Ui���c/��uF�� TH�oI��>�(�  ��j��<�9�]P�����~�ڞ�n7b���S�� ����(��'�v�Y_��:�Q5j+ʤ�*���A�{�{ɣ~�4� �f�l��}�JX�72�=��Dϵi�V��䋖�����T�^:)V��!{�-$�D�Ь�A�����<�Y�-���q�C�?{������.l�2X$���ւ&���%��Ȭf�t�g��y�S��3u��}/�-\���Ni#��X�<���i���W,&R���֨��]��n�Q+�v��g2"|o���N89��M$�+�]���)4 �!�G�$����G��)�g��Y`-y8��c6r���� ��ǒ��UɆ[P���{&�y��������"a�]"�ͤC���}�"�I�B#���?����ii�.Mq���3=�'����6
�U	M��d��\��pG4!���ܚ�ЛRu#q̹�Z7�<VA���`m�;�o��_��jDr	����'�Ӗ4Q�	9�-z[Ⱦg]�˺
��:5f���uƋ��,[�L��Y93B�4��3�
/\����}��:�X��p@���	�C�$c������.�f����qY�&)$㈏ҙV�$ر�6͆�h�\O)Mk*\����K��b+�Y�כ�6�R�B��9O3K���#1
�c���zp�����tw�q���w��*��	�r&�����?����(�)9f���kd�ևT#:���?�������F&b�7E4�Vw�ν����a^B.�e�Ud��)A��� ���-�~C�K $2����Ubq�Zk<�����
�)#��zV�ٷaNץ�*@��B=bs\��(=��곌�ˎ^.�#Yg��g���vB�.b �v�������D��'(x����{B���*��!.3Dq[ե���О�=�u���ʿ&�P�c�!
�C%�2���KD����@!w"ðHTv�>�����<��?.��=����O&��BӸ��U��y���=D�9CR�u
��o�n��t�0�����㷖��Bid�l�&8k���!��2�����#؆6�T1��2ĂKd~�0c�Jgo���z�ʋ\ Қ�|z��e�P�dV�QG���Q�c�6aj�L ,���n��L��|����-����yz��nB�U�ƕ0q{�p���s��W6m�[w�x�a�U���`v��A�E�"s1�����&x
��M�o
���U�ŉ�Q�P�
I��q�Vz�f�����{���4-,{71*�>��Qf�k�|�mq���y"�N�ㄎK%����(�������(�װ��Ԍ�*��hYp[Ϫ).�tq�'9`����.�'-j�Kl.5���T��b�{�r�N��t d�
C��J�87�JR���J/}��Mb�k}�q��t���&��C�g���BXQnܛM4du��P�p,�2���1�8!f���c�� Zt��pq<䀱�T-��Le�:��w��~!��,F;�GS�k��!\�io����3����D�or�K(�|o'2�+�\xգ�
4#�ا|��4f�(�ؖi�l�茮.��<h� ޸��Y+{rX[��O�<�ￛO�n#Rp-���