XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Z�\����Qg�������{OP�X�K83���n�Ѯ�~}y}�R�\2�)뽀B.��Q_B+_&�����$��يG��#�}Q�d�ܛ;x�/6�7	#�Hdۮ��3�՛�K@y؂®a�|��B>����Qz���E=��{��3���2��qyE�ͬP[<*�@<��I���u��ԭ�N�ݪwXS�l.���>.ИƋ��M+d5	��[	5oN��6�*��p:�0�?�솴|g�F�f=��m��e1<�ly�c(����?SeL�"ъ�N1F�p��rc�m�W6:���R�ҳ+�<q��o2fU���AQ�,ۍA{%��nn� �!�!ı��S 2��D��5�|����Ng��t�Sx&��C�
XA�p�'�'/�Y���ma�Y���t�zґ���y7�W6�I݁�(�p�{�+��p5����g��a�c��`�$����M��Z�����9�n�ҹ��v��k�c��@q�{>��cs�p	,�HI�Q="�=�����+ˀŞf�� �9"�T�+�ꨭ���ݩ��m��^{?i�f�G�	~L���݉k'?������TX�ۖ��Zc��wz*�����(���C��㽈�!.�8_���8�%%p��p4q��F�쀦gr?���Z��#噌an2M-ӎ�O��@g�򱓧9炦6��5O��A$�M
��#$A]I������U�����?Y>*G�<��ޮ�Ti>�v! ��@�(XlxVHYEB    3fdc    1160n�/��+���ɑm�s����7�J'�`�/j�4m��(R���-.��~.�P�b��u�9�=�8�m?k�l���a�a�ד�E����N4ԙB�Oȑ�6l,^*x�Y�g�?�%2CQ7p��d��lP��NA�����E���1w��3��=�D�p%�X���hu��Bz+��Z<�0�� 	Z�zh!�J�p�&&�����ESY�?�#��(�,92���>�GP��J G���GO��9�I���aۼ���p8-��tv���N:�g��׊�	�n�^���(;�t�o�,�׳AF7�^�4?��0�t9�h8Ԏ��h�����7g�<1 0��=��Ki���Y����}|�B�^W%��c�(1#2���a���S��=�;�k#+��E�QKRP�;�����{���P0>O�`��AՒd���=v,�
S�F;vO?�F�����N�%Skd�0�y�7�
����M��ԛ ����/M�E>�O�QB��rT�2�^�/��C%/9�-��8Һ���Ʈ*/�9x�/ҵ��fe��2�t
_�l���ߔ��K٣�>�J��v�Bu���:ʔ�E�����~�o�e�3ndkR��߮�a�(e�.�L�:?����K��*�/򗆛AZ�q����p�f �΃�`�ޗ���5ckE Q�sAmN}
��V��M�j
V�SBs�ԡy��@����Xʲ>���$D�i���؏�_;��W`˧AK���Ob�K���gS���"^p��@}��q�_�N6�I<�AU��,�w��ŌyoW�0;؊���Ȗ-�!����Q��M'���'���Yמ��1�T�c:|�$2�Ĺ˽�683O�<��F��{��uzﷳ����a�$1ņc���2���Y�	��hg���-��<������pUi�fµ�5�d?]���(�a�n=���(iq��&]��	��bg������%Z��tM��>�4h�M�G�4ı�N�t��k���T��N��U:��ژ��'��#�}$� #~:y��g���Y��E�b:#�N<�wCO�Xp�S��.fg��+"�-���x�ʔ�|�o�������a�����n9�֥�o�G�{D��^cMt>�� I���5�G�9�{� +6�)��7ڢ�Y�E��ff�ix3z_X}�"��eA��`ytBu�.Z����C���e����}ϓ�!p;���R!�I�08O�q�NmKF��Vc~e{���C�VaF %\�j��)1�{c�X#����1�y��M��6�7���dL�j}D��x6[y	�k���U\�2�3��ZG� �_N�b�O�k�sf�-f(�<���w{'I�ݖ�-ɬ��:?	�G�҄Q���+>M�H�SZ{��	��l7Z���p���!O=�_����)%h��@��AVI��@��1 ��ϰ�DqG��~�惻ئ��w���Q�vu��R���Y*�+E��3�r5ê�a��hٱ��T��;*X~W@(���ˈ��y!c��1�?��bO�I�
�=��dS=Y~VwY��I]�ރ�#�Qy�G������H�q����1>O	�����O ��kw^���.���uzF�K�KC�� �:�2�Ѕ�	�@_d����z	�oqX}�~�l�9o���B���؄k�ĜYς �XT}��Ju9K��/�-�u?߹I9a��%��y�>�A��k��-=0lR���b܂�L"�pM=\�G&�ڬ�x-��]P��eE��[H���C����q�ɏr��ܝ �i1�i�V)ʨ�g$��2t��ж)�����;=� �)
@�#
�����̣�C��ak����A�,���"��@�;Q�ff3���aH7	T��F׭p��8�9ϚLw�vW5P�WB�l�+��͞% %#e�׹��`�>����Y
5�\ߴ�E��B6F�G~�% ����_S���RP�'yN�j�'r��s�l�0�O�1�"�pqK�Ɯ�uݜi��h��t���D���U5�d9PX���H3n�3��u�(��Ha S�-�~�o���S������AӦ~��IE��4��2ݮ���#-�fߕ�^�T7�:�vP�o�qg,y~1���R�yE�<SK,,&�6���[�f�o��m���GTew��k&��9�Lut%�C@.�p�vE�o�3�0e��>�͹�~E�,ZLU]�� ce������D�N uZ��At� �}�+��k^��F*���T�-�9 4:­v�FPr�>,$���"�5���Mb?�/�K֖H�+����b]nL�� ��-�!U�հ�.��w��$�i�;�����R�Z�I�R�6�Xw��+���=�l�*Lj��a�e�<��Tsv�ي����Br��Hu,5�P��u���)�;Gx�, �@��> tuP�+ô��ϱPb�ڋE�觶���WҶ�%E<�:!��3+!����*׍���E������z���/�){ۢ�
�s���Y���8�&XE��Cl��u1RF��ׄQ�AV&�ӌjo]�3@�u�z��8�W�_�{-+�O�g:��?�zR!�2�Z��W����3�u��Jz`<�=`�!X�K1]` ��d��0��N�FAp��3:�xrh�Y��B�QzDp�p��������wl��=��V�}�4�W�H}8u�Q��.�)��10F������k \~�%�B���b}Ј;���q����W���*K�n��dT.tV�Q�hT#f��a+��ɗh�L�pCٔ�=�G:��Rϊs��[s]�Zxs�
8ww�a=��z�آ��4D�d=S��.C̵:*���m��8��뫓z�tZ����CX+�=�b�0�ac���8䣀^\�
��0��-<���J��,�*�Y�e��ɎXvǟ=�d2��o"�vg������w�o9!�g6P���[��JK��
c���r�c��ᾕ6r\�������5L��v�?�� ��� eX�x{o�������/�p�Iۈ�fD�_��8��ʛ%>ۉ��-��"TYj���UGF���mJ֓�ދ�_V�Τ�<�^�+l�7E�X���f�
���Y��uش;g�T;9%�#ȴD����%�;:f�z@vҝ��iR�S��ź�W�n_���8���U��u��+��:���k7dejժfbѸ���t$Z Vz{���i0�?V�`!��V���+22u��
#j$��t�ޫ<H��;�#�`b�7�~����<��O�Q�`�1gK3�y����
�������ɸ9��?3͆���CM�`�vYp������׻��ijtfޏ/�0AP�/U��$��߶n�Wo�F�|�	��x���)���]�\��S�⯷���&���(�n�{��I$���جE�㐠B�ُ�I=J�I��ۜ��֎g���K�P�ɑ�tޟK�w�1�8h�}[�:�[1̯#al�j��(�u�R��D?hu/�����0�ڏ�d[v%lI����	�#�I��_��V���&�N���JSK�pcӍP.n��o���[=5�i�ա9;�d�.1M���^�� .Cy\&�*AG���my_���qo���/�%���Vt���y�%�~��@��R �JC�ڜ5M��I���E)��:��s0t�����xO�y�9��D�=��tH�>���c�<�ţ�)4�4'�a�CY?�#�=Bv�}(7���������I8\,���;�ˣ�lH����lS&���%�78^V����t<�%[�&B�9F�����Ӿ�Iu��Y׌N"DiL��.2K
w%��ટa�<�C 	��
:Eԁ��噢�II-��Gy��R���:�	�@
�zt+��u[:!�xG�M{�
��	J@��I$:�a�i3;�q�Dkk��μ�I(`L�3�9��x�۟���	4[��j���g�I�T|��],:�n���:Gl0:�h~b�-��yw��)�s:-g˘��͟!l��%2�]��� P E���R��5�Y\`�1��������:�kļb�b��G^���K}���;/�m#�4W�h}^��*ɫ��/�Zh3/�H�)�Od�L�_�`̳6�Yb�OH���*�գ	�E8	}����l��޾*�K�2�	:BO�jǐ��Ԇ#c���NA�nr:	�[^�]M>�M�(5!����Z�W��`Z�����)z��u�ڶ7��%ݷn<�Vs����)L$�`8����O�����i�c�.��Eugkr��[i��&H�'��d|`���	U��>��5K�u�
���i�j�[�l$����H�Q��Zfo�Om��_C�M�$������P��ږ�᧠�T[j�'=�qjx���9.��鵃�~PK^������Yk�mN��n�40?��,������Ā[J�ˢ�U��c_�\�mJ٩ t�3�"���0H;I¨{����+uWM6�X+�tW