XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���_	-t0�|9ޢ�pH8���4�T��;{m����
����ż�d�ߥ�O���y��c�֑,�\�����vP��ŃWA��i�Xt_���@$���z���ۑ����xoC�tG/�DK/�w�0�4猜?T������"��G�}�'�s��N/���_���о�U�V�[ɡV��Ρq��x>�`:g��� E
�e*�cv�{���1(�� �ۖ���z�)[�|�N�І=#��,����X�FO���n;�����#�N'm��
��c*g�ݟ�ֳ�k�iMGL��y\9��z5'�,���y���ʪ\'P���e�b'}G_��@����]l-I ����o�b}�TrZ�G�h�x�"TJ���@���n�")D���r�Z�Z�P�?�dE�d��uNS�f������cj��Ѧ2@_�t���4��ވT�Zb�VZ�j�Pk��Y�M9�D�̛󈛛鲳�㉓��=S0c�Ɵ
R�5�����Ҝ����������`4��z�a,L<��������0�u4�4u���>���?3�����!�ǗҫS�h�y���8�-~g�5YM����QZ~��q��u�Ą��ŭ{G-\3硄�.�z�JNx�Ѓ���m��H牣�C{��8���B�8m,_h*E���s�h�ES���	#bOG��M�*!6Z��z���|�s.�8b:�<AM&!F�!��Ug9�X�Uf��\2�a��>-��*�w�N�e���72�Y���XlxVHYEB    42ae    1110�Ad0#��djf�(�@nn�O�~]�r��~�/-�9��`��_��A���z)�y�r��/w��|�+�Ps[�.�̣#�q�_K��[K����j>*L��w��!��\�t�A	�n�:ȯlov��)X����R�lCF����ל*��N����Ӽ5#��|-���w�4���n�&m%k4���'�^�{n�?=8��"D��^�|�u�Ѱ�j�L�]c
q���o�m�8���0�j9�H��:�@8­7p���tq��㫦�[^~���.Ʒt�!Bc�*�Υ�v �Y�T����9��X�m�p��$E�K���^��l{.	k�ABg�!<gߚ�#9��x��2�X�cӖ�f��,[�B����'�X���iI�4�1�%���i�`�K ݻjY��׎BOH��|�l����Հ+����̱m�����ύ��{�ȷ�n�h���gspq���n�j�!�#��Y�����}�4ǆ��ӏx2��2H�9��e5Ej
}J�5����ѼUhci���0%T�~/oӻ�QYJ���ȍ��4�n��n��<V�*�l&��ѹHa?����T$�ŧs��ǎ�2�iųm/ρ�[�+���I�ğ5FA/ggf8�!���ѱ�Q��pb��};��H��A��D,$��W��J+
�<:�7!�xJiZ��Wj`P�~�n�x�}8�����:�����zy��W�M��_��ccO*,�����WiU#����-M[�)�b���&��/��6���Q�g�>5�1�̀�H�>K�rh8��^�B�e����'L5�&"�B�r�9��	�)~�6$����xp�SqM�7�PT�r��u}wP�"�-�|��v������������M�����-L�P�N{ ���G�s��o��34s�w������:��J��!>R���<���D1xK"� �cu5�	���7ꦞ�����5�o�W>u�����کh�w` �l�����U{�/'�~)�&�� k�:?r���x��\aψ<�H�V�~U�r󁒻+�Ϋ�ms�+BG�p���K��ԣ~d�2��h���.������閱r���h��f���+,���yWg6$�!����:νe64���Pʫ�s��n���1|�;��zP;`aj�/ka�#�@/�������V� �&�0+�k���|X�38��.`!����C�W��3�{�o�:S�#���?tf�ZjQ�ށ����勃=�vΚ�i�I�U�y��~���[�_/;��L��FӮ�4���c0�Ic�P"�-�8C`#<Ʋ��&�a�F+����i�Ƿ���godi/@E��О�ҷTT��bރ5�G�_����/�8����񩤯űX'[6�U����ĥj��:/n���3�!��}R�z�T��ъ��,�^�;n��:ؙ�g�����*���rm�h����?�͝x��trC���)^m�*ui,�cG}C8�C5���9��	��?`�m�bW��A�K�r���Vi��w�:�A>25��Cf5�t�ȹ�,���E�w�E�������F�6W�
Bʩ�1"='3��(R�ƈBSZ�@�7p!ݬ>�EF6�n�l ~���cw�|vYҼ`��GF�Zt�BQ!������_�(㑡C��n<]�f�R�T5�t^ڼ�����2x�������(�*<�++I��� Z�[����E6ZV	k��R�eT?�-'ii팤d� %ו}�uZ�m�G�@M���&���r�����L�H�����)����$�}�ֆx�8S�".�#�Z�l�qM �3$�[K��m�Cu��&鞑s�E�ݎ�bż��FK4/,�;F�����H(��;�`�U�*�?+��[���~E�b+�	Z����Z�6i��+�F��W#��FH:~��p)���Ys�)o�3�W�����-�/�Cď�ҽ@�`$�u�k-�X��ci}�-zr���)��y?���?ŗt�y���Ɋ&B�p��,�w6�ڀ �{G�9~R%�Te&>�#��XpJ#�|��.ZhǰԤ����!�ߏgt'L�	���K\����e^��L�t툾W��=,��g�+&y�tJns���N��F=�p�}^:M���ev��n��'O�tl�6�7V�#[5$I�H3����~�|/���l�|f�Jö�o��b;]B�B�r{��k��n^1s�@�#��f`:x!�tI>����c�l�Y�>Yp6̓��v��z���qJ��m�8��XIVP����A4�R��E��+'�	S�&ǽIY]��Z���0ϒ���3�n��� �KyT=is^`"ml;�1�5è�m<�"��8�se}��ˮ'��n��S,/a�>�aV���&�IL���)���Tc�3�P�<6w�g��dT��z��"/W��~nL؄%�rH�@�����]9ٺ���.��E�}	1��4���g��O9p��P��%g�O�p�- �ܕ����0�2x�>�����R����QH�R��<���У��l�r2�����W��-1�P��VYq/z�g�R�t����v����V{m�d}���\zFէ>w�	�H%����3�t�nV��|�X ���zyZ��f��q78�pt��h���#aw�U�ۡ��̩8�[د�P�
 ֳ�#J�u���Й�t5�x���>¢�����`vt��T^����B�����,E���ONMV� �G]�N��>��8�dU��NB�0u�շ,̩�5e��(��'}f���Jp�}@���q�]�
˹��׷��@2��5�����b�R%�Za(.����~5[G�ǵ�R����װ8bV_1*���j�D �	Br3���Cs�_���q����������Ud��@4J�џ��=@������_l>��2^p}�$�7<ݪ);ʓ�`�W��Z�q&O�X7��g2B<�E��n�"�r��,@@��m��Y8�r]�m�A��K^uz<N�.��H~�T �d1���$�ϔ�S�:�#���'5Ս���_��Nk��H,W������f,@6&	}[���d�m�xPWo.�$�S>Y�X�}H��-I"�e]�Y�?	=������rO�H���ro<�f��fE˧oFz���}�7�m�Y=�����Y�aF��<���ɉw�8���0���O!P�}��;�4&�KP:N���o�t��t]�a�Oϐ�U���±=,~0p����G���r���m��4\�&w��Bv8�@��!� G�"\�r�j`6������@r�ԛ6��kIy�=-B�c!��ɹe�B�nN3��c�A��U�pF�s�3�o��ʶ�x��.7J��%��*�ѧEU��r���C�٧�43�gX�y��С8p/z�G
�PH��}ܸ;�p�9�&�h����#�)4��Y4���ے�r�͔����aI�5�5k+�k�n�7�P{�	���}��[�k��#\�!�g�W90=�b����u�E"u��$oAd3Ii�ml9��3jD�75��$l��X/��T4MbO�kfȺ��C�<y�����G]�`_�lV\�a%�T�N�n�S�.����UMe9TْF7�P#գ ��ǸQ?ק���/���ۺu�4P���o��l ��o�_BMO��.�1E�%'h�}��-z= ����q��|0��Ȑ�[�K#�/�q�`1婅�'���U�4��S���޶�?^V��s�&z��I~�9 �#�ԙ3^C�t�k�������u{Dn����(����Wۯ� A�G4�	�>���PGY�华ó�:}
���&���6�)SX�$CxN{8�8G/U�f_�@W�fM%,�)���C�=��l�b�x�j?D�C�zK�HKh�hۅ�p+�w�V����eCQv܆=��*t���QV��*�H3E�����)��͛� �����Q]��I�F��{�t� �J��Y�4C�<�܄���V;�?.���%��cʾݰ�,�}�p
�/��+*�i�\����9�z���q�He`�E��B_7�]�ۃC�(��������rN�){W�ϭ-@O財�W�Xe�_�ް�zW�!��`R
�r /{�*�A��~=z��kAJa������۫��w5�-7t)��S����XAX�j�����c@��\@Ϣ�	}2�bc� �����,��70b=���b�=�#,?'Zz�Ρ�*D�积�&�4V^��%��ڬ�00	���?<���_�J���&Ɨ�PԵ~>����eV���U��A�Zʜ]�i�m$es�Y�a��b2�K��P^!n�Em�8�a��ۗ҃�a=�N��Ԙ