XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��d��V⌞'[��������w����
!���q�x1��l,��ѻ±���vQ���v3��Vz.S(g�
�x]�ϊ5�Wo �L�$=䲈*$�p���>�7߰�����X�ww�)�R�$���N�1c>͋�ŧ�]��6h���B��X�v9ɢ��PԌ� p�BZ�S�[�����X�aS8߫��a~۪������%�Ȩ����T��Q�=6{>����OF��\�s�����t��}�.�e���m�*����-X#�
����u>�I/�L�/!��їa:�Z��h��v���S�c���d���̿I���S{��H��f��e�1���ʘ�l���4}	�N����#�N�r��YMVTȋ�
��"C׊��:�d�Qq/��Ϸ�|a7�C���.̂H���b#����з]���^W�����~7Ɯ����z��)m*%'��Ȉ]z���� ���~<�
�h����hi>����6�����%֥e�)����?�C���?�G�܄HOr��ZP#�������ԉ�C�����H7�;R|ϸ��z��g�7���@P�X�l�Ի���Η�ko�����> �s�݃�W�ɷ��{h{�r�#�}�8�T�疭.R�����b�ߴ���U�a������r7Z(����ȃ)�H-��I��~G�ީ~���\�83\ٕT��H���3}��=ިA�����o��br�%/=�(�d�.��T�H�WCXlxVHYEB    6014    1840�a�����_�Ŀ�pg��h�'L�̗��ň�'@��h�b�.��X����/�e�Q�(�!��/�� ��{q.��G���0@�!+=���S!\�.�f�=l?^׭���DcG�#��W��J�v�6���F�%�M���B_��
 \���7�a��d�;���JX"�y��$lB�b�5�����]����v����P�W�3Nּ
V�>�֠V׵�����U����8`jU����*4~���$��H�7l�����v��E{i�kzD��>yd�ͪ.B��h��XT��`cw�&"u#��=��M���,K=W��^��K���-O��t�(J��F$� Ʒ����)ÄQ����-C�7z�A0������a����� ��O�E/%;�8�VZ���C�1�^iюI�6��Q@A��	0<r�"R�Mq�b�Z��������>._��QB��,��W�os=EJ�U.z1Z���cuu��I�˘Y	s��e�)<,
��C�+��6D�'uo��h��;�$��Hij�TIA1�*�:GfH>����eh�˻�ӠOƌy��eI�.6��^��c{<G��a�@�:�2����w�Q:����t���`;ϸRO#�7Y?�)|�NVm�Ŕ�Ժ�m�����M��GE��6�J�]U�oi�W�����3s	�w�`8M��K�'p��j	'�Uf'���ɵD����s��`� r�0�F��Jx6�M���9�C�[}�41��6�Z �a_�/�����ꚣ2}?����$���Gez�{㧟i�%�ۺ���{Ę:�$&���˱#[m�ԋ�%��G��?(g���x�v^,܎��7��!-Sx�W19i��T����.�+�X�eYRA�H�@Q`7�Lg��ѽ�'VL����:E���"�����L�L}�@G��*������s�Z��J�"�{�gQrkt�o���� �n|������#�A.Zz�� ෾q��nPM��BU�rLZ ��_�Yy3{*h��S_��� 6���f�/�Ü,�h�VU��
��Pv�8�~�+�E���'�Ƙ��� c#���N�)R�I:t�8n��]�D��f��R	#�P�&���*�FQ��v��|[#�� �d�H�O���C�c���Ɩy�f�3��o-����S�LuX��)�p�̇� ����3g�\d_����赊qbq�S���5�߅i{d���h������B��@ƌ�{�Oѳ�(A�������戅�5}6���,��$:�ơ���b#{J�O��c5�)6�]ڷs[gH�!P4w�&��[|�-�;M.����2�մ�>�i�s��,6�g�ȃw]."w�كZp��'�=P���Lk#�G]�<���m��{d���
h���_��c�Yy\�k�ٴWB'Ht�AT�B"�'��ʺ
�Rdv�-*�臄ÙvVq=��+֩^$��&NKKB���� ��g�|����I��=Ѹ E��#/�#�9�DC˞��{?�.|vc�Gm���8�0�����wn�h�b���$?�N3��n��yW��(���s�'TR�,�_un�$�xk�S�nF�ZFVS/�<x2�j�wf������O���K1bK�L���6s�{f���BN	 ���#>��!�eb�Sm��k�ュ����G�%��t
s����}�����l��t#�/����(��\��邪7J���J�uΏ)σ�B�
䯣n�C�FF!SK!�.OA�B��m��,:sۯӴg���U�CvAZ���d�et3&��p����T#�FA��m�sS%`�oA�U�� �{�q��M3Z�����U
H�w�-[�"�����ǹ�<=�e�u��,��YE�� ]���ê��w��\q��Sh���vp����p���9�r8��ЃSy�/�YA����
�_�'G�p���F7���{j��t���g�����~��*��T��>B쫊�N*��~0�����
�!1T�P�f��w�Wg����4d���3_������c���}��`M�Փޓ�����nW�Y�����҉�m\}���Y2�Ѐ���;�I�KB?�_�l�n����-��>"��q���mX؋�o��0Bx�)!�y$icVZ�"�w&���e�ӎ�|���Ǝ��/Ԕ�b�e�Q�L0�(�պ��L�H��Ƚ�ڈ���;fx�7N�!�nY��ݮ�rP��k���^�\�.�E��"twq�v-ˋe������;u�j�e(/�:uQ�{ܴ:���h��Mu��<�����[D�>j�
�B��g���'Ȇu�f>�R�8|Z���ԣ?�����q�$d���[�g&b�3�V���S�u�U�����ro*"x���C�L*ҽ�Ռ0�9t�/���;���f0D������*H�������ƙy.-����̐	�٢�~G��K\�9��	��&��Yl�&*!<���?���_�e��֏�)["�Pr\�4&v�L�����0J���EvMd��B������h��L�#��	5��A�0�$�eq{p�)4A���3NnoD�c�S�m�@Ⱥ�߉�<l}+@��.���s���Ө������$w�l�6�����U���b_�8Dy����[Ŧ��amrPM�o��*o��IK�ĭ6ۂ\���u4Qp�A2�ܖ��u~�ʼ9_�`0M���~z=��O���wĺ�jvr��;]���VP�SoK�]�MPƪ��܋�.���?��1���+���dg3�m��%݌!va�̒��K�K�k��-��"7���Qc��}�?�a���(n��1�x����X���%��Zb�/�`.�c���Fq�1��:U$x�<P�Zk编x�}+�<��br�K|ؕ�ͬJ���)`F�-{  ����q 0����9`�J�b[���r2�w��PsF'sT���(�h�I��@���/��TV>���G{�- ��`�Zr7�p'_���Z5Ƴ'����lS���=��	�E DNQ;�WD ��=<�������v{�[���P!Kqt�d��_��%1�ܷ��&�E����'����g�S^�B��I4!�@��"�!x�=�ŒP�ϵ�wZ=�WPl�l<���~Hv�w:t��6�HQ9\�f�e�b�/������ܼ-3.��Fs��d~ �2jqt��{�~~[x�֙>D���rd�vh�@���D�w�P���%�F1�/W�R��Y�̱�*��I�xR��N}p z��ϋ�H1�C������Z�^�\kL�udr����0�O��6�}�
���¿_�����d�D�֥|-H_�-�?��K����'ʎN߾��6+[Z=����\ϯyˢ�~��r�p�����2݊���������Z�w�^���iSb	��uD�yH�<,���&���mT�{��'ҏ��f�˞��E���ߌ[i-��-mu��D����)���4�k�>�П�ӵf���fu������S���?�a~�)p�qD�"g�OK�$��c�f�L���:��!���[���)(��g��ǭ�Ua��y����U|�h��u`N������I�� w~N�?J��fM���௣T��A GR�Lq]�:>$���
M�2fve�̳�Y~:���'�jrC:d��u�F}�������T�3�>&;%2 �9Kd��Mk2[�l1P�L�$�B�4���(����̂��(��x�N'��CM��;KP��m�'�� ��|L-�K��`w��m{�~��0��nB�[�N#�_���)G�����cN�r�?z/ΐM��.��o���S\Z�>Cr1ő��%��.m5��"�Q��$C��aU�N�a��&9��6Mn�@<�Q��l,��B��o�*iN{�ֈ�7���;�!��CKM7� �R��;��`����x,��D�n�C9��}���7�p��>�[w'��u ��
Z7	-��"�a����)����! ����d5z�ں���ϝ(Xv��){pt����yzW�Y�]���`��AQ��U�e��4�~��s)Q�'%�g�*#�Ч��r��.��<��Φ��47�	d�!2؞�b���./L���=�Ul(�x��m'�݉2�)=|]���G2�H3�,����F�#I���G��_g��Rc���c�4� �&&�����#\��W�B�~�ؖ2i��|�ݿ9���`Я���G&c���y٫�He BĂY)�� )o�R-�f2'�,Ӷ��Oi�(>}RCv:�n=YۀnG���1����~j7�*� ��Z���qW7�
�n���V���m	���lvu�X
���-��{������5�neI_|[��f�A�-�e.�0MU������9�8��N�����cu�*�p�������\@e[���ڡ�zHw@|��X�ͬ�E>z�8�hW�R��SR S���	U5��&z��h�㆟8<>Dn���qA�{��{����oPG��≳V5�=�%��p�����;�AOch��R��yE�@�',�j�0p��ο�݃��U�?�&l�ڼ؏i��n�S��"8�-�!�5�Y%
E���A���嵏�/I����Xu8
 t�eP��`P�@8à4�:�uݞ�>�I� |��x���|�}�LV(��'��{�e_ĵ>}N1���u�E������#�� }d�Bervt��j@���4h�/8�� =_ꗬi���^��+���?
�2�_�q�ǅ<pq����N@�2Y;ή�4Do�L���E,��W6&�Ôw�b��ѪI�;�a��$�����$�C+~q�4cy�))�S��@ǉ(��x�Bj�;�0p��׏��}�Bز�^`&#c���E���#-7�������-��_0*�H4t�����@o���%3%"�sK��kƷ3�{���f$�W�]�3�L��j�~��1��|�B�2z�c0��P�k��^�-�R�+E�A�&�fL��.'ţt =�����jT���5�Q�*��fJ8Uf�FiYY�Cj8�J�´�kyf{_,�k�K�4���[��i��L�i��d��׫rE���k�o��8`�MgΦ�EZ���Ju�1(��۰��3����FC���O�?@���V��t�.�=�UxNoV��H����=���-�Q6��j�Ei�2$��]c�����u{喩
=�h�D�LH�f�GKa��pazç��^���E.q�Z�\���Jp/E*�⋤���"%���m޹��~yj�4eJ�8{��=P�-p'i�n��#����+l���N1���oL����n��	n��7�T��*��(�l�MC�ּ���v(��wo�}���M�ZpF�Ʒ�A�n5�X��G���D�P�$�y>&=|�N��H�g
Y���V���۲d�{�gu"Ƕy���/��2��*�tf�7�����̀�@?����D�:�M���#�DD��d�*�]���񌂆��4�}���0�"_r�4`z7��؀֦/�7�Ă֞1�sK��c;�@�����E����$
}�bC�|A̡Y磑&g��u��ㆊ,WL���l:5���7�d~�$�H��н�z������l^��8=����RYE���r�^R
�~򴦰�������ۊ�4�d�ӼeR��Q��z�G�	����{�p�/���[纯�/X?
�N��N��C�z~K?�����=ÖU�jK��̵�3�f��6uq���s��]�k����`O&9���7Š�o�F�8T�l�(zj~�-QӠ{i9�#�Lҋot��S5���Z.Sj'���Ĉ-M�l[�bs���n5��[�2Acu=s����^�I�D_H��|]�U�G�7��=���+a��#ػV8Yde[Ł��ϝ�ݷq�}�U�Fq�K_J��R^���ON���Vq`��z�K�?#af�!��3��������]zN$@Zg��ڄ�}�V~���g���̣8�j�� ��Z��_8��4km���������I%O�9U("�\&{Htl22mt��������`��AjH��U��T�RW�HI>�d u0���)��e��
��3���`S��
��P>bo��e�s,�