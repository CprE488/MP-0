XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K����� ��ab��\� ���K�D9�<L�� �h+Y���Y�H���;����S�b�"�7��A	Ξ�)i���V��.������n߿��]��ºG��N��^�I����爀�t��;����E0@�-3��)4AJ��4����z$oo5���w\�yC3�G�^��h���o��ap�η��m8%��Q,����5���N��W�fN�c��R�]V�oA�j�2^]��l6����+[��T��/qp��Q�p�T3��u3C��f���܃����}��h-�lA�-L�=�oL�8�7��:t�e�2����d�'�ZJ���Tٱ��� ��ʳ�`9�<+]�,Lv<<��U6.�Z4>4�fB��0��+�L�F�,�\a�7�"��ًaH�����C�� �A�]��q�h��.��V�_�ֻxw��T��%���و)����"������u��C: �wk۬�tBi�u��v����sk$\��-U7M��RÅzA�f'�1!���f�7��Q���Y!�:�c�O�=bF��%��߭K&���ȝ}����͖��͘��wz&ӿ���I:+�*L��l{�L��k�?�Y�3���
_K_�: �ng������ʠ	5���O�#Q�U�T�iO�.ae��}�&@`"|ȨW�2|��f�G���a����(���N=�G=�����Z���F���O���z-�y ��Zc��������e�r AqP�$�z�@�]
����z�XlxVHYEB    6346    1790�t���P���� }�� o�y�~�ńHh��M\�����+.��^��']!q���xfY��A#73CW�wV`�cZ�}Ц�����uY�"Y�$ַx�8!��Y��$��nn|�qc� �-Y�ڻ�	����a&S(|���dȜ:r��ˬ����5Y��X�F+JA�RY�~,	�i�y����\�W�:eK�2���aZ=�� ]Y�;뤛JJ;�qF!Dp�jCxRFLX�ڛ��w4�$�KC��Q5���t�(%)��wM�q�g4.�&
�X�i�W(Wd;k��9��{�[4�����z�}��E)\���R݃�`S��X[��ۭ�7��cg|�8��H��\| jV�mZv.�/|>�U�)Y2"Z�>=�HE�����.lh��3'��J9	��们��e]e�xG��e�'���pmT{Z��)t�}fl��ڄ��]x8��':�󙰀\��ݶ'� X�B��`�Ԡ�*��|��KԨ��8+`�xx._�7��բ^��0���X ߞPY�)���:	��X (�b���y���t\�dv�__�}�t�D�L���8�U{p�,K�ޡ�N�X	�e�$sw	ܯ� a�w��p;�]Q�5����Ta|�+q�Ƿ�#��*Cc��[�@Xբ�wk����"�>gDZǣ�����S��� H�t7S�#�+(�Ո�[	HLf(����1~�@(
�Bm��W=Y��z����`f�1n��#O"�T9��I�4 �R��`���k?ؚ�R�K��p��>�3[D=�|I�8t�7�V���*��T�g�7 �{��R��-1uI���.�޴��p�|�S �����<��n�i� S:�x!�g�k�yk*���J�92�u]� �w��Rsx��*uѽ�\�� ��N!!\��-�qO�N�!��lh Jb�l�/�wh0��7c�����ћ#>	�&��?�!�$�%~��n,n�\���.�U���eN�%4�����R>�p�;Na�b�  ��Z�ish��A�:K�x `@��oqPa��?ŌJB��?e�Gw4ɏ�Y���{���"�5ǵ�m�k� ;#��\Ԫ3��v)�I�����&�g[�kU�W*��c��mi�C�(�P8*0�a��+J��|}]�1Tc��3����t�y��1a�|��z�Bi�Z��h�߬	s����֓#���-��O 7歓l�!Iaܘ8��h�g	 K�9�f�GM�B��#�T����U���lI�f�"����[m&�by�SwU�#�A�tC�L���u3�{�����DA��qR	��Tڷ�h���8��$v������5g�,�p���r�/Fk�h�*�l�:�"%3�Ua=E	��q�B�'�ԜޒW|� l_�׆S8[DL�NlPee�s˛U>��a��#�P�I�t:�16b��7}m'^�k�_�%�k��f���ڧk�T��(�?��f��<�H�������f�߅U�=�#��1	ȮRu@�ω�!�h"������'�ɯ���ak���N�-�JqXw\^h�"h�E{rR�7�a,�*B�e;	����b۰'?Gi�T3K��ǉ�p�AH�<���ѭpv<�'n��^��V?یd�_� ��y����M�$ĕ�֤向���Zl��ޛ���t~3,�50�g6A��Y�Y�����XL�Z��9�O��TtUٵ�'�=�d6��n����>7t��_r��o}�8����2�0^Ɩt�/ޜ�p�(�k���'�O,�ox�hp����i2F�?�T��@I���/W�>�p��}�Q�-Yz�ધN��� �QU;G�RB��j�Ĕ��i�c{��\�+m���d{xIA�VI��b�AQ�&D2�]Hr��D���/#wԿ[(�G�uy��Z7&v��WD����2�{� ��p�*����g�]TgހX��:s�'�<������X��w�^)�3�o}U��+�յS�kܸ��lf�Y����mq�̃{)���-�/�w^���餽!Ԍ��:�hڗ����x:����
�����ђ�dl��3�mQ��&mS���ϣ���O��\�BS{z���g���J�G�]�-���56��Y��|��e�b�8+z틘W>b���<o�RU��k�,�K̽��	*�9A~'e�`Lk�R���[U<�b��� ��ۆ��:i%�v�aI��=xiH����
=$���K{���c���L��hjLV����0����X��l��;��q��E��8
�4�C V)&<���Vi5�ݬM����lf}?z�"����ƔZ��6����e5@��ڌ�C�e쁚:�!�5�J%��S��5��V mU���؛7�L
�*��(��7��V�S,e���0>���W�L�Ȉ+��ih08��ޢ1G�J�w
����B��XJ�T��C��7�թ����:�19)3.�>�>����a���E��җiU��f�ɰf�ۄ���p{�	�1x
����q������˛�� ���i�ˍ�����i�&�M�WY���H��/��
\�P5�)oy>%~K�B�q[�朗�`kݏ��a�ᙱ�G�����}�y�3� ���+�Y�&{�f,'�"Ns�=B��B�I߫�b��w�z������Op
v6�GV�{	%����?z��y�|�?��Iݗ&��D�4՗��m��
����m{��!'�
:�p H��8ImZ��aa�}ݣ����j*�5�L�rpR_2-�Ř�0h�����̴���cU����qA~|����!����8�#X��2����G��e�o����h/��T�4�/�\d*w�f����>���$>��co�J��E���Ŀw!z�N:���9�4g��� M�!�p~�49�R����*�!�%0cKyP�:r���v�����!|�Y�9Q_%
Q���!Ɍ�|�+k�wI9rq�4�� ��B��u��ͥ�,%�tN�AS��61u�ZS��e,vtiX��������{�z��� ���+��o��Tq@ ��"��h��y=�F��k���)#8eɯ�T{ޫҰX��ℭˋ�_�76�d������Z�P�.����r��i�J�pi1�+Z`I'r}䞙�C���<����5}uhD��o�d�g�X�
e�3s�M� �K���,��Ad&��RU0�_��i�����~+f�C����x�>��^��b�H���>�ۉ�Z�m��]/%U8��/̗��^��&1H����ՙ�>z�fa��VZHkG��P����t������C(�X�M�Z����#�D��Ǆ��UsY�_��i�e�6����c}]h.(��d=��<S��RC_ �;�2ϞO��<�6�R����f���ʼT�~�M�����삨jV���ڳ-�4X������X�t�
��f��G�{HP��O)A1���2ġ�0ȵ�Y��<OT-��o��y8*_R+��K�y\�/f(�nN,�@S%�GFзT�0�tH��ܩ,ƭ<�X�9�30r6X���]�;��6�aAi3��ܱF��v���Ѷ���P1ɾ� �*� �%v���hl���R�Cr��ȿ���_�2��t<u"�`.%H��k0�����J11爫��ބ|c���ƽ4
/5��uč���vʴ��S+�뻮�F$���6s���7[?Ib�}-P�����w�`0T�h��%�v�u$�4��ƿ?�{ʡ\�B�bmĠ�H�\`X1�ф� [@�}��\���N/K}Jo�������X"(���mn-j�v�g�/F^����Y�4�{$	�>��
���ԣ��:�J��������?8)hFa���lA�8�7f�x����_�k�|�4)����v�_GXX�K�����>m���{#=r�~��]�c�~D b��Gd�� ���GQiIFҰ�j=�+����&��
��.�p@l�b��3PR�Qh�ߡ��;�Tv��&}DF��v�� �+�������&ln��D���v2�^HҭI��h{{J&g���Ԕ^�P���l�&�yLRE��SPb+�5d���j�߿�ʐ.7�T���H)��<�����嘙���h���^/�\KLz�m&�q�9�G4��h3� �Bxb%Qq�X����ί�@K�9�LEp��N][�S3��`��*�<�̓�Vi��U�Tm	6\*{O��i�H��p �o�5�d�v�N#�w@�n7'����D�P��Ia��c<N�����q\�0�S���G�zwK����-�!�m�f �w�:�Y˨��(�/��nc_��tHa',�b&{aƆ�ʸQ��Er�7����K66��N�O�u4UⲐ�8c��K<����mz��觠�-��3����f;���{{8�-�<���x��p�
�n���5i�O��Sj��54	Y�0Z9	�RhT��r��O���(v�lFј"��v��/�o�Y�n�9D�d��$ �k��8R
h��4�slO�@Wz�L�yk����<���6eO�[��?��#��������p!��0PuK�����F��x�z��/�����r��s5W���K�t��A�������t��YwQ�\��e�˹-����a��`��B+�1������;��íqeI-��"��{	l����"�=4v����(����:�v���+ћ(�\�T>nk8���4�_�hp�%^�zӋ�I�����`E�.��;� R��T�茝N�O��t)o���a�}��)ҙ��N[.n�u�;5����Xv�܆�F�`��L�Z��8�^ȗ;~�W�V���!�iۇ��Z$� �`,n�-(�w�(�P~Ւ1Rim�,�&'�Do�&���t�la�q�I�Cb�᧾��C���ox�����G`�L�	&�C��xv�k�`D5�ˏ�i��+J ��E-��Vh�����5}gv��
��3��ic������K{X����0�s��U������[@�$���-p��x��=+QTq�?�D V�?ubƬ�����e'�[��l#fJ&�?,Y��&���î�Z������H�
�g�
t��ָ�>�-���2����:��v��0Z�s������ |���=�����1eT�D-I鄳�L>7,�OZ�Ϟ�ל�P��Oݡ�7:1>X�Z������V�C^��䙒���?
��=t�H?�:���X�y.�K�S�nh��T��r��o%�.mi��C���x�E���<�:�TI7 MPE��?� y'r@y-�Bs����H�W���z9�����!�˒x^g|c�87阿=�Á~υ*��Zy�7_iUB_j(t\�.��+�(Wɇ(k��0��Z����Qy��&g�J��Y���i�K���]�_v�ڝ��
�B�"�$�U͈���L��wY����Qި�xb[p:S;b��%@A�4�-�|���/❼����rc���e~L�&����'�U���g4'g�(�u9��h`�	U\��&��G����;��HA�\��sӘ���%��m�pdx��Q+��Z�`c�E2V�׸g��O-ۉh�آH�L�s�aOiJwV�Ȗ.������μ����f�˨E�M<A��L��"���Vk�q���O�s���}|��n/mkz�!��ʹcTo�N�Ƭ�m&oZ��B|�Y��m̤N��4�'�tZôI4��nRG�>�}��z*g(���*��H<��"��5���@W|�ӑ���)�j�Б����,��3ͭ��͙�^_Z�3c��k)���ʭ�wJc�ޏ�u��g2U�k�<������#;����w*�)�WYl������9����`�`����8SN]��8��Fɗ�R�jm���*��ʶ�d��r�jn�[�vT�e�D��M��"-\)E�|�BIDB��{����u����x�L��"b��,�<Hp��$$�n�I�9)�e.y�^PO)N^����