XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/{�\�V9-"��%@rs__��C�- ����Y�O�	Zn� �W((��uH/�,�Oi׍^J���QV��l�3��@]lD]�gt52-t��9:���7%˘j?�g���"�z���hje�]^�{���b$t3[K�s�O4��i8�)t,[�l 5�4�� @gST;H�;��0����!ta�@%�/;��b1�� z�,ֺ¡�7߰.frNĄ�4��l�����7v��j ũ;͈���{8N��?ح�:o�-d8�$Zl]���s�L��;|@���n%'~}�Aw���?�W*gX���&(�9���D!M-�.YrV�� �f� .Z��cZ��t0��J�9{��S�9	�a{a��\��vqL�#{:kQ&�� �]�-����t��i �T���SvF.u�'�?6cڭ�(Uh�U����{(�I�k��<?�h'�<�� ��g|Gk�_�|�Q!�D�/�P�����=m���v�#k�yQ�|������g�)�RCe���WT�s�IU���4�f���n?�+ z}C��r�N}��ΘP�j��*�ʝd��V�dsK���'q���gj���� �tS܅�8���NЃS�Vf6X�u��#��+|�G�%��әl|rȊ��>gE�f�J�0�� g`�~5"m�ɔ����Z�y,�Vo-��.���n<�~��n�f�n��2��0��&tD�L0�u�R9�������3"O�m��ya��)pq��t�:~.)�F�)mXlxVHYEB    95d3    18d0��F��o���ȟ� �	���C�����Xh����k#I��}u8��jk�܍J��	���OfgZ�x(�h�+;^�=�8�anj�ꭶ"?(�x��)V��0��x�7�g|ٶ������|�*V��B� *1��ef���뜙��UǺu�~�q�e�׽c}�Н�
=�p����ޭ��!�=����\��Ί���Ο��/�7BvK.~���� �n�C�ԋ���/h*w�
9���a� rԅ�&j� ;��:���LNZ("~=�U�]	N�Ʃ)s`�e�cfY`g�ŵ�g��O�F�/�HR�;�����ɘ8�&�	b�V����d��M�]0^\B���D��!�Έ�`���	�W��Lŕ�r|��ryt��y�b0흒�4( ��q "{��<h���3My��a��8C?��u�b���@��/*C���r:{�kj���b�6�#�rp��]���1�����zfy���b/(�T�9�W��]g��w�1�"���v ����K+�y���}�ϲ�`Sw'hx�s�eLb���-���r��(&���5�����_�mW��P�u���:U���oߎ�I�_��=���D<l��վ�T��-m��ڮ}��M��l,`	�x~�ݯoF��>÷���݁Q%J��8�7��lC�b���QE)�i����$f:�Gj ϟF���P*��Aj6� lN3�&o��+EI!v����cgP���z�9z�8| ����Z��Zy�����K����B^��:�����q����53n] �[[�k�5# ɳ�o��ћ����LG��q��G�`�q�8�B�U;ļ�+���]�-�X:�&J)��qu��u�eh�]~V��(�mai�.��2��ȑ؞��{SBi�ƣ��2�8�Y�e��Kʮ׋~�ҙ�t�y��ٸPcz�l�G���9�1e'�KI��⊤|(UM��N���i�|���F+kKv@��Lbz��hWVb�%���*��4��9[��A#HOH���%Q�LIo�� *B,q2kw�����ćf�޷wc��Q�0;]�=�L
��}D4�+�bC�L���3.�ֶE!�Ō�JJ%3[�LW��xH�#�;�����x?�}L,p���wG<`���6U�M�e�v�Q�+�64@�\nf>�}Ȓ�.6�C8�*IM4 ����~�8%�1c�@�#8���,�V�zA}���#��ʾ>��G�J�(��Lf�I����f�N&�ny4��֥3΋K�ӍW����Fr�j��	D��>����o�2�6j����3u-�_����nj�V��S�7�� A2�Je�v�2�j$r���T=i%I��K�2��V��e��P~_7��!	�Sܡ`��#t�@wd�D�t2��S
<M�������;I�w# �T���؂��^@���dKp��o���aT�RG�A�k"�6K�fLe�I�/Zw%<K~��S���ܶi�ޕvщL_Y'	m^3��]��E�����sDW!� n�[���6 � ��i>�m	��	=if0�w������ą�c����VQ$�P=�\�F�Ф'���T�0�biz&�J9Q���u2d<��ǫ r����r�Ż(�����.���?�mN��t�n��ʫ�̈uU���%��������M���Gn�M�.P����{{˒bXA�u����
8��u���a.[�Ŋ�
��5nL}T�
��kN�an �Q"���^�����zf�V�Bơ-�wm��7�,��t�������K���eS�TZ8t#���c/�8��/���sY=rYKI��oK���׃@t �JQn�u;]=B�j��@���wOS!��g��L�"��f�/!D��}��� �Ó��^NV�p�N�Bg�\Nt� �}/v����:0�#7d�C8�a��5$�E�I:�� ׽qSM��%BM8��Zq�5�����J�"�G�2ɸ�Ό�@�X�U�F�D�r�C?��ĳ�"5(���}���u�dn2U��mf��8�X!�������VN�L!��s�`���X�y�H�nZ�]h�XZ����Z1y�j�ՈB���(0��}"	����(u��⎉��o�<���.:���gz���DV��n%���&�;ɭ�l�7��l��D0hLɊa>&Qu�`��1��	UW��ٴ=?`i� ML�Qkh�|��-eht>���6��5�%g����lⷳ�3�L~����gq$h��ri/��J��J?�hI��ɚ��BG��n(�2�;���e��f�-@��m����%���u��G&�#����u��U΋��=��P�:�O)�-k�\�=�����Fٚ[��7G�e3����ݳ��c��U��Ӛ�CUG�" �N�jZ�������q�\u�8��;�b��p3�,�h��?��p�#��.��W�W�[t} �6䦅���f�/nMCr��H�Y�7�"or��x���N;��zM���<i՟ځ�M�?2q�x�\g9{OH�=?��9D4�IEg���:Kl���O-����Ϊ#׹0=	+w7��t>�[��^uٰ�_z��>�R����͍�?m{wș�D��.�H�C7;`:I�'�E}�{bdD�!�c�\��t���Ts�Ռ���R8¤����y�dЎD�滽�e�\V���٭� �TM(zN�w_W�D&`��
�>�,_�>�֣Fɰ��*��	p;��̍*M�g���WZ3"��#�^���ݟ�A�Ku"�k�E2�.[�jB�GAG�W,W���#��V���Tf�Z�c���j��bQt*|�(�0Z��SX���s=�S��[����l";?,0+�567���$QwT0�h%� 8M.즟�Fh�Tݢ��z��K��^�%~�` 1��n�Uْ��IaM�"�1QvMf}�NfE����8�0�6�Z�}�ٕg;bZ�S���>-gBmP��ɴ��ŀEKE��[�*�F��k0Z�-jCd���gH�w���q��e�}X�⋩�#Ru��^y�C�����O�P���� ��a<��C'0@#A�C]���Cq���%6A��A�*��iOY(u�P"�	�hJ\b>oy�K�М���'C��f��7n��"J�E<2�q���B�#���G(jV ��x�
<�D8���\@�;5p�q�J�ɍ`e24�J�p��4m�I�g���)��{��V'n�V��\W����w ��s	7	�`�Mt���VN�G�󶬑\{����]	�[��|ue7LJe΃�L��;�L˪�f Y��ʧ��������i�R �]�ӳ��[�;�&�{>4v�#�Ĕ{�t˷���݄=���>]�E���%1��zpL<�L	��Y44��kZ�s��2����k�kT�I��Y� ��-����k�o�uF�6N �"°=��f3�e�mE�;������h��aS0���u;'t&�}<�I�X�DК��Z���A�#Lӂ�EWL���!n� �~�).�6��`�vs�!��؟o�4� 7�'Z��+Y1G��w��%d�~�#�,B皋7jN�{���W��`��#�/���!�������u����+���2޾��vW��73~d�;G����42�,��F^k���Tx҆��p�G������r�/��l^��(����G����� �ExJ�n�#�~3�1ҳ%v��@��<��Q� .�E��5�YA��h(�?�o(�+:��B��C�����f(�>��T�j�t��=�܁��|b�n�@
�CG�'��,��j����Fb^o��oz��p��C5ݟ����x�+	-�n��B+���~/���b�Q�*Uub��_j��Zxc����� �{��9N�Q0���:f���ޝS���s�?��![=\�Re�䐅=��t�Kmx����(?l�b˻ۈl������ZS����Z� �`����_��%�&��0�����:%��0DHϗO�V�굀0�b��g��j	R�S��})�x(�.8*U{ي�8k�D��!s�DCԷ�d�3`�V�#8%�-x�������ˢ�0���w��0~?� :i=��)!�lB`����E� >�'��4 ��&�ř�}-�@�;�ODd���%��a����%&��մ�0LBX#�P�ypi�[KI���������(H�7����Ŋ�!�Y�f�0Ei���U���|�7�!!���d���|����:V�7˿���H��L�'���j
g�bK6��
IcR�L���t�,�VȚ
9p�=a��_�Xı�*�8P�Ԥ���U��2s�-�~1Vo��R�9�U�]��s����t9�ŦCg�����Mj8g�r7Y�%���%8-豾r�u�K\�f8�Ԡ�̆��FH	$�X�2>D��
ϓ���%�\BhXnp�wfu���=��O�ˣo3j6t6T�t�rq9]㿕IR��o7L��HG}\}���PPka���)������pC%J��Bi�f���{�(;���p�c�9x��n�����-�r��$Lu�z�Yi ����"�����}���4x]�2#��nȓ)J��m�U�ut�%*�0Yޥ���PϹ�s,�
��K���Y�b���#P�������Nt!��k�[�"}�^)�,�s��)�R�w
t?k����.�߯Mf�q�CW��hZ�R)4�!&סڌU�+�4kud��;�X�2:���ӽ�R&Q�K��],^t��qD'6��$���F٨��K2�^�N��f7�"�i�{5��v�J��?�dh�<t�d�N��?	<^3���#�Ĵ�
����e��(��� 2[jF�g�5���+�ؓ��.[�I��Sn�e9��g�����۫=� ��xU���wI7����;�X,X����O�Ǩpl4�e�ӭV�Bg�e'�^ՙZ_M�HM���83O	389��4iM�K�a�ۇ˥\���c�8�fp(�M¨���z2��WGN�	��s�+/�h�?�u�M�3�ke?}x>� �9>_���R+S�3�Gw=��ҝ��B���4��4m��L�|h[��O��� !+������I���?(ma���`��{���zIcG�=y`q��X�iA��rh��c�;f�n�~;������jA��ke�О��}w2#�/п�,��Q�'.�1��	kzkw���B��E�e^#C'/�׾�k5����-��#���6m��7��'ַ��F�]  y�����M�7�x�Q,u�U����/w�Vv����>����d߾�t�P%�?���~��eC�9�ə�M�+��R=c��7qa�P��)m������@����-nE;���!��X��0���v�`fj��M�}R���v�����.]RCR���w���~��e	��
j.�Q�2ӘZ����r���M�cZ�#�n�{��D�bY�o��Hy���5�d��5��J�%g�L-��7�.s?#�gGBZ�<�� /{<�פ���l�����k(��ʸ��T�ש8�� :���2��/��b�F�|��_�L8Iah*($󹕏�C7N��=�d����h�G{2Ln�V�M�E�Tds��y�uI��T�~7�'�G�$^B���
֞O愜?Q7����֡�HF@핱Gm鹜ò���۞ǚq��x	���G�qr
���B���� ��
b�٭��8j �=���n��d��}GF�|�#pC��^/�9�:/\H́[�o��HD���',Dd'���>�Nn��$�(>]������:���^�7Ae��qo�����>N±�����è0��qaѷm�R6*WT���L�گ8��nN[r�C��J�
4�E�F��Q`>K�1�U+�|8�R��
[�$;q�d�u4%:_rة@ZT|5���UҊ��~�av5������޵��+)�������}3�^h��{�-5��"�Y��^�O���ֻ}��U����G�k��#�)��kZx��Mo�.�u7�1a�R�ǔ����Ð��2��|{Oe�J�ð)2�kQ�SH���/�`�q��X��?eg��p�O�����GᲔ�0T:�Nc���b<ޫ���qp�nQAJ3�UW���4�n���a���ej� 	g (�G��*LV���}�ȫ�%�O��;f~d!�\�ᡗTј L��D�>f��6������¿��'���[$�S���m��J#�7k�&��8A�Z���>�r�~��ŵ|