XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G*Srb>տ�©kz�`�~Q�����!��&pvA�هbV�I}:��\*Pj��$���q���!����zyn�0'{I�a?U��5�I� �h0Y�{L'&�:j0f�v=�)�0�9�u���+��j�ӫ~�� �"������d���SE=�i�[���~�2_�oz����)!W���d.z�8���0���M������o�ߝ���-OP�Q@)�@_¯[[û��@��f#��T���K�w!o��L�4K��s��r�g,�{��G�ڈCt�ۨk;�O��Li}�Y�6=kVSʹl]n���>0W@b��e=Y7s��{?���,*��e��:�E�ݦ!S�179Ӫ�~����q�VG��Z�������#�O�&� ����ˑW�=XM�{�w�Y��k�x�<�.g�+��[��[�J���-����SY�NJ�b	k������@P����eX+A��UO~������%t�Έ�	,3�}DT0H�-�H)��d�U:q���'9�U�}nF'N�PS\���P�)p�Ue�Xw�A�3��N���5�Ӆ�͵ '�	�*��,�3�8�Ү���\�R�$���*�/�R�j�:G���H�Vc�je��ۑ� e}u�ũ:r!�r�׮���8�Ļ*��Q�cN��w)���٭�uqwK��7۶:geȇ���S������$�[� W�e�}��H���l���1�v�<؞R{�C9N��& �8��f�tXlxVHYEB    6014    1840�P ��X�ؿK�b}���F0�ʏb���/Kp�b=� �ќ�A�0h\60� ߗ���MOs�].'ߖh��D���ά�y�(QŜk�(�e15i�� �W�YVh����hJ�Ĳ�Ou����
z�h!�7r3~��'f3﴿ƶWo���
���6�@n�Ifc3��e���h��%�>�vdDr�0�"	���0���(��CP6�} D��]*��e>����TB{
g��a�ZbݹE)��h3��[��I�x�ERֻ�'�5��`S%0b�#��º����Q��f��.Hہ���X��ǧ�`]��8:Q���w�WJ�D�
6��x@i)�B?�L��U:e�Y�����Jy���gW+Q&=Z+���8�8,4�<����3x�J�1�J��u�|C=�xgCỳ\	bb����~za'����̀�c��R9���_L�(���T�@[s��9�����Կ����܃t���#W��O�o�?b����]L5%��)Db	�[���i��=oN>�5��tF�v��;о��d��=�RF&�?@E����k���S/`���`�8�cPR-9��3|y�е�b,�di{�����l+�^~��c	�o�+zJ�k0�2��)��
5�8��šizT�@|#��
t6xgB}N�ZⲺ�~���Va6�y��09
�4�r���Y����2(/c��)�i���	�� Q|)`=��\x�;�.2�3�8�r�wC�<GL� Y�J��Ͼ�)M'�>ٹ�Kuy�" Q:�T� �Op����lD��D]�R���X��G��,ܫT>�ڕ��N}�a�#p����"��6�I�#�W���1Ѽ�b����%f��͎!ڱ_��q:�Q%K�";5��ld���&\�������讣��/L]1�*Ċ��ԏ 6�z3�=�"��VA[=���TOy\-��4�w�9�ls��QӞ�Y$C�u�f�=�W��׿�J�!"#���p�����mNm|�kR$�&ޯX��l^����շUpG%]W<�H�p�TA3Rk�|q�J�s���Ѹ�v�t<�&[��]�$����v���O��� ���<-�Iɺ�"9Ɛ��],�Hfx���ht;*)t�������N�1�=8�M�0 Av�f�d��N��,����2��WW"S�DkaP{���cUj��n����k��GyC�ӡ�(�gܶ��,��B*�\�4��͙ ʿ[���؎ǬeJ-��Oߴ��џ\0>\U�������֜����"q5��@:j�������ɖ�U�}*P,2�=�I��n2�`HSۂM�]����$�,��R���D�u�����.Wja�¸�[��̧�8���B`3��ⱐ���}k�כ	;4g��37�5X�oD	{�ľ���8����Ƴ���	J͍|gWn��lbr϶&߲��k���|�M�O��U,�;�䔫BS|VҞ#LQ�jZ?��L��t��b��S�ڸ4�2c�B��肕��fS�=ŚX�#N;6������B�\ �[�@�vdR
�� � ֡ӗ{M��˹
�����Q���	�`��Јs5WG���	Hi���_���	��F\c7�*����0��)	O�'��nܕ_+L��6�"@���r�Iyl�Ł�4��[�ᾡ�����1�yݺw�[ @�3T������j� Z�u��(kcmt-����b�-���s!�N�p�IFgD5�쨓+!�����~3TK���}5�!=v��°�R$��aM��+�{a�$(�Og���O�n�A�ː�	yH:W���'B�bΕ�m|yl��
}�.�a<|[6U}t��0����~l"��ӲH��Y����)�H_|g���J�c������HՄX ղB���zQj�����O,O�oZ���%�!���j!��(F��+PWYȁ�E��6��Lf��Kv�
z3s�"�#&l��4=օ^
v�m�pRu5E]�j�?�~OGЎ�6«����c5�;�A�
?l���@8f\�мOS����;�>;Uw�lI�#e�׭c���W-�H��޼+��<hC��O`�!�HyUs���?���B�����3�{T,��׿���z�N�T�$H�Cm[�z�K5�X��a�j�<�=���E4�v�(����Ѝ�:�Ŝ�h�,��8��XH�����^�W7��5�E�ׇ6���e�	 �����'�fN\�Ʌ��Q5C��	�	�|c�_Ա��0�	F�+2�X����7��U��¼M��b^ۆ7���|�Tw��Q���êE+p��6w�����(��T����efY��-�F4ppo>��H��du� �wNk�4 �:ߝޓ/噿(���jSN_�H���~m�Q��w��ճ���A�':�v�!�ѕ:���L���
#30\5�XE�si��)���b;��C��� ��?U�R}F���P8�%��\�QV��*`_@d�\�d���G�HEve���,�H4���e_ŋx+	H官��v���Si��C	z80-w#]�����v�U��ɵZk����<���Մ\b��:��G"���ᧁ�M�6\����y�A^�5�����:�H/�s�
(�߱÷.���!QʂD*��KCfhҭ���p�!�E%��٫�e`Q�bu��,�m�n��O�ٛ���qÈ��� <v8�[̬��A���w�������Y�g���A�h��Yv#ճ��tr���m���k�q麁�������A����DE�cgPW%By�������m�v�x]<���@g�9uyp�NR^�Y�_����V�@���;}t��ow8P�1������y�e3!�Hr�#��K�L�S���!9��I���c�|��5��ˈ�E1�DN
ѵ��e��%a`���w�Ə~H*����`�kQhHan��@ % ��=����}4>0BȧQ������6���	K��
��@��f��T��;��R��
:c/`�76BQu������W<��WC����.��y2u�*>��ع�=�����Hg'FT�x��^��U�����HM>�)SUW>}��C��U8�y��^&G��N.�zr�\O��noSC����9�����W?�omqr����Z%��'���M6Apa����3,f�A{K��Q�ȍ��m���I��M�"�Dc�5�M���d5_��i�2�4"��p�x��~Y����.h��!(��Ӷ�����TPe2������Vt<���q��C<*�0��:�d��S�S!jK�V7���u~A�Q�z��cH�u���./�T��v[㙈�C��~�\�	t��
(Gm�T,a	,Y8��+ϑ�����߁K���|1��sa>��@qz��yI����>Ja���!i�Do��#��v^�͡gk���Ա�\� ![��u�����!ƯxX����3�6���}F	9Ϸ04�t���~�9��\S���,HqO/`RPa��!W�m�rLU3�j��4<�ށ4`Ko�ID�E�˭�K�.��RU��V1oԱq��7Q�5ͯ�(K iiu`Q�pt�q%�L��Ԟrd��%����~�X��2���|����άE+�]�1�|�����s�Wo�9�=̅c#փtQ��=�RԚ�*�b�2h����.��!�%����S��#�$�)d�+��cIi9aI�?�yRM��o�ôF�&��Uf����~]=K���Ƃ�M��<e��,����2`cFu�J�ѯ�L�� ����Ֆ2q�y�t��'��s����T����	.�<�r�N����{:6=�j���DO�q=(���53M�Ѡ�\W��*z������Lj�X�J�\G
+Q`h�L���O�.�2�XWƿ���q��jY�ػ�����<���&nLV!R�����"e#��0(N�G�@�f7\� ����Je�D���T�<����^�uga-m��8������޺��Hm������K�8{ߜ���.;�b2�_�ی��)%�W�g\,�� {;�"_�Ԍ1A��_fE7�*=q�|��Ejr%)����;��w\�`���:'�Q�3aW�|�Wg/����x=&#<�؈��/�H-a�'knd0*x�]Č���^�d?�&�˱k� 
��i�O��i*�����s^<q��Զ� =|������|���*�0hyT 6�w@�QA�xp��4*X��%�b����I�ьiI\�%�P�sSq���a����8D���9��J�,��R'+ʹy��]:)���C�VxU��Y>�C{�?����=i�F�O��/L�5*��p�nx�P��[Hm;��.�]�,ͷ/|6�ջ"T�gy�ol��.��>��10�/${�(- S+%�B�����u�-��W�DAk�,j[T��|'�[��kҝ"o�"]�_�P�����w����T�6�;�0�/E<�fI��P���i�oF�P��C=��u	�P�'�n?'��l;�F��ݡ���M�b��M�Z�,�`i���~�X2���'��a�����Tg7�js����a�즘���XM$��Ӹ�t�������v
�'�:�6�bxDan��p�s7�%�L��
XH�E�s�9��?����h��pC���_�]	V��Զ���Ʌ2�_���}:/�T!���[r��Y�*������f����z�:�
:�!�=p({�˱>ܚ�gF����%�*�V��i~2�<➣h:a��i���e�N���>��=�ŕh�Ü�jm�
��J�����i,��n�� ���No7`�'v3_=a������&�(��K}`��|z�q�]N)�#1�Cjɭ���n�_T�a�1�����â��Q֪W��%�Bd��y�<%��͌!��vL�\&<�J�5e(k��VF̵y��%����5���<aŨZ��+^�k��Bl��� ����,YfbŸ��*I��#N=n�T�Cj1?8�U��w@(M]�E�Y,qr�ڨpF���@����#-:�a�#u:��R)0��M���	V���P�-�ȴ��`��xf�~�� R�:�R�1G��N�)F`P�ɤz>=S���\�d5�&��E�}��fQ[�2��+WӴۋde
���[9�e�~e�{l��o<J� P6�3eSQ��6XU��FN{�h�>Դ �;v'9y��6u�}iK�^DJ�&�.<^)�E�� ��0?Q�慘��핕�t�K���fe�������!�� ��)�~��}�`�����+l>z�DϚ̤�N���m>�o���a36�����e�F���A�SqmG��)u:��q�sp����kB+^d�o�]���]J�߂�7S�55w ��gh'��=~,KsG��l�v��W�pX�>S,���<˄aD5��%	}'j��0�S�]▴K�V�1ޤ%MLΤ����B�G��T��Uರ�o:MP�� �ٝ�3u-2��e�$�A{Te���቗c**P�t�?6J��`���a)��BuN�~�ih19A��gYF�Mn_C���}`�i[v�S���]�P����\�uA�/�Y�����A�H��Q�*��Q֠O8��B�}����2�\����zϳ�]~��T�U�wzh9^�	��w2��MUH���9�5���hH��X?7�~�.���;O~��o������S�\�rQ�����P)p��J�=za��^�
kä��5�J�R�"�o�"(�T�*�.Z�D��0�e����S��߂||:*:������שԝ�z2������	�rU��0�-#D�2� =�U��"7�݆�X6��(�!l	�[e_O ��h��Y��Ug��	��?�rMN��q�����W�W�os�Q��^)dL�=C�&�n�F���v\�1�����bJ{�C@��b�-���<�ۉ)�_j���3h��*Ỹ^i�V��}L� �����\}h�d{�;�u�A��-��	tV��NM�}\�sm��BCWO�!ɷ=!��Y�u 4�t�Pm>�#?9�����|��CB*�q���L}�`��/����I�_����pJ��w�+���U��ë?��5=@
�SDz&����)��_�-�s6YP