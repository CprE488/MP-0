XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���d�C�&]D;��.0s₩�r��7�qd�fFY�����)�ĭ���*Sȯ1�C�=|K�l%ZT8��H��3J/C�_5��X|��8��&�0}��knd��Wx������fJ�r�Ps@8���<FX�G��!�e?���{���������
�����\ED�<����OY�]�@xAsbA�s���'�߽�^�(x:�q�GE�Οkg/�'����%E�`����W��>��g��)Q��1{J����z�f񙊤L��^˪��H���n ŚCQ�(���q<TL�?�B	2q���I��Q��7$�b|����H<k��4�A>��p�GǤ�B�x��|�D�����L╻$�)?]AG�T�>m��z���=������#�Nl��׶�n�#��4�=�+U���%wNǙ��<ˌ�Ϙ☃j�l�:k��"���.���(�>�\��]�J�m�$�m�"+/�ϑ|i����8W���rX˻W��E���~'O~�q3[]��)�𣭲_ؙ&8����j�6�a�xm�X�<`��)iG�O�����>D]�n�[���j�up7 �䋒�1�D*T�=�J�|���飗�<�i�����X����)�|��E-�e��j�z$���^<��Jg���:g�Q2���_X����=�,��Nv�x�~�y�]�(��I�k���/�Ł�����*�Č��Vgj�$�V��G��{ �����,<�+o�� %�[�XlxVHYEB    a037    1fe0�K�-i���	�zXsffB_���E�%���
ܸz�_�w�jR�|$/åV�@�Ov��)����\E��.����H|c}�F�ɞ,��0��V��p��I|���O
��^ ��l�$5�@��r���F���hu9}��U�[�!]��+nP�o�u��G�`�m��M�o�g���U��طS����nK ���?k�,�p��R3ߐ��փ�Qg1fi����Y~�Ƭ�n�Y0-�7E�:&QW^V0t�b�7,�_�7��_&k���EHخ4�$R98w0���g�'V=`�|]��ǰB�A�Өi�/�Sh�b3.	#�Q|*P,%�ႚ0E�"n�a	f�89ED��t�#�1-g��4�FӢ���+�Ͻe:²��!#�YlY�m�0�O,(\�d�!@�l�~kg˙P���KU���%
��d�(ц؀�z#��~1��>)�&��E|��6��x+L�k�+B�A�\'��0�L��E}���i�-�D,������~��+��K����m, �o�ZR�c�[ƍV;r� �B�M�%I�z2%r0)����{W�p&s��.�H_�#z�V|JQ 3�F;5����C���Lҷo$7�*!ȣ~�<i��m�%,j�� �3g��ʹ֥L���#a��z?�
|$prFW�rg�ϊǱ�&	h����`�q6�s|0Bu�#? $��b��W�����b�V��6Q����&��L�wGb���T7l�#bQ�L��;5iΙ!�]���1&n~^"�4޹IEr�.����iK�8����[�@��{�_��������$���\��P�XϕS�ɐܽ���m�?G�*e�kNW���V���z��[v,Hf&=���zB�Tp�swd��b!�S��7�z�y�HzK��h�]�0~s����� Vl����w������B�a���P��T�3w���]��S���ZS�;�#�ںS�CF����q���K�J�(�VX��n��M�o�WÛ� �r�ܷ�����Q������>�s�#.+�o��"D�w�(t0ΣH�8Dm���.�$���Ig��A���	�xk��`�/�M{-UY!���VWa�|;�6s�ӥ�i��EF�9$r��"c3�T欮�Zט%	ק7�m�����n�۴����jyU!N�Az�6p[�,���i��Y;�r�$�k˔�L�y��FŌ�t �BM�V��_�D�Ӯ!��p��@��[�~��D 4(���C�Y8�%Wb���t�c�g7s���9邧����0�,��CW!�\v�v�j�3<��NGD�,�?n#G�`u��5��EMs�@�]�u�)�.�x�Q�2y��8B`p�[!j��[v�n�
�6�^���U�"����֫RmN�u�.���=�Ѕ$��3f�dE��.�M��-UX�l%��l5�q֌U����U@>�F0F�+��0�TD�Yh/�I�0�!π�O�=M�_�N2F�8S@�����6'�i�x��\c���4�Z?Ԏr�[P��0���-���um�G�AG�q���M�lȡ9(yf�����r���2�����TV�LF����N"����Y���� #��'�2p�O����`q��P�-;0�����҅�$u$�[���m�<R�u�;#��#���ӟ��A`l�����w����q;ǩ�S��ڪ�� ���"�mN>�/�BJ���4���(o��dWr>c������}�r��zd����o�3��������ʜ����{ˏY���1�D�ޱz���@�Y���'T�!Еߴ
���װpiu�"
�h�;6��G�0��Ysm"0�$�jq) �Ǒi$L���y�A5��R^vz���b��Ic�����6/�7d�q��'@�nӾʝ]�o��%����J��P����;?�� ĲU;R�*�5��8�������| ��~Z�oE�0��k�c���i�G�Һ�h�2M�@+�Z�ui���IT�j�	|����Q�[�*QY�*G���,���@I���\}��)	�!t�t��(�@���k��D�4_�?N�V��툁WtJb��yq%�gkc�����e�'ƪwv��L��I��i���ڞ��7���z�^�y���Z���< v���D�E?}�������~��L�ݿ��J^�в|���;ē��xhU]���F�R|uK[����E�^��͛ F��JwnL�v�.+D6�?�q��w��onk�R��2�J�T�N���N��A9�N_4Re���y7	� ��<١�"V{��Ȏ�;��͸.�%�B\+Mj����2E^@iy���Gm����g���v��n�- 1��lӢ��|qW������w����p�������!`)/%����V8K�b`&������d��r8�BhuE(��rk��	��=��	pd#Y�t�3���qE��my�C��|A��sC��?PK�,�N�$kӮ�Y�#k!S�6��f%�(+֏��Vb|���#���酁^��_o���I����gd����S�02�S������Wl���_��/����KPtXK��ϐ=�!�w�,�B��Ysp����S����c���.�>�\#�Me9Ȫ%��dXmX�줤zeL������`!5��<�+Κ�icA\A���Y�ej��I��blm��\��z���ņ�LB_��qL�$��v�354*�(�Y�UBR>X���=i�4�	"��>�
�ػ|�8��J	i�J[tzL�"[8��r#\�y����xs�ݦ�z7��ϋ_�R-B���VN<��pƳ#!F���4{��V���R�"=u�]�E��=.��{�!*2X���g�Ӑ��%6>)�T��yv�ַq^�,��G�f��QW>d׋�����+���g8�&���T��M���L	3�� ����41%��-_xO���W��<��.Ǆ�n:��^�Cm�b��1������lPӦ�F�~s�F-6�^��*�/�����JPݶ<׫+���^jv��a���?e��4�!�]D��z�_�� �eʰg��0�J ���UD�t�io�~Q�V_6�T�F1T���7�Oϖ&�;��o����ޘ�'�F_`Z�%�w{Q]xT���"s��9sH3z M׼�ɂ-q��޺��!�O,�c�N� ad��~����ʊ�����*A�B�Mv�7'�Di�*6���J�j�FbK�������?��I�'�n��k�-e��g{%�#Mv��nG� \���ϖ�.�b)��D�M�z]��g5hO�����N�`���Ԭ,��(o����j��b�xD�Z��ܫ���Pe����s��m5Y�>�*Dgh�h��� ���p�8��~����tB�I�����ɼ$2�'���&�3�~��ځ�#��r�����*�i5[4���x	A��AOB~
%%uUO��̑���pi�G��Jǹ�Ђ��	����%:�z)�dLA�mt�Yÿ`,��6F�!b��L�a�,E�]%sk��+s�z�܄�a�OI9*=a਺�Mg�_4�4��j����k��%T��+E~Lc�����Y5:1�m�v}Q�8�K���s��Id�,_D�v����4V+�]��vǛ� ���U��q�7\UU����j>a+0g$��A�a��*���83Rš'�@�N�6�85ʹ�D߸U���(���;��H���tn{3��iN>���N�z)���|I5\��I�gW�� ���KKx�nSl�N	��!�G�����)>%5q��A(�P����R�B��PDt��j�o�N���i��$�vL�f|�����E��M{��Y$���l�3�������t�h�2��uV/O�u��-�L>�Y��l�ѹ��Y����֩��n�����B"�A�����Pa����Y�j��|!�sjc�*�!�3���]E��j�<t)ıɃ�-:!^������7}�����G��2<��5W+0ڍ*!1T����Nlo�*B ��G���e��f�Z*�V�E=)��X��e�2�WW�w�T^�,�L�I�wq�	�CC� ���d�~s+��߬h%]���ahz$���[-������B5�M���g_�
Q�}�\�R3�,���d���NÏ�'��ff�Te��L�"�lw���9'D9�t���4\c��Bnt��i�u���@1��8�x��}��L���T���w4�ڹɠY:�Fo�Z����
��N��(E��e��6��O������q�2h��m�	|a83�Y�*������Zx���p����b��E�Ok��}H=`�^�u�!^�:P�8�n�i�-N2���l�`��x,v��	���.l{��;O�Zl�4��Ae�쿚wn�y55 O	�}����k?_U��0�JqP�`P8z�k��>j�gˑv51�����"yؗ�[9�*���*�)��+WV$���e�1/��=H����VX�D"��s�i
!Wkߤd8PP>�?"�Z����1��~#�0�4N�Q�m)�1��/��A�'��TR�;�8���'�����'�f�(Te��}���m�t�w6���q����eeF�[0����{Dupa�4���A�H��<L%�BV�Ym�p��	�6K�L�u��?�� �ӔY؀{�5���F.�͝u�2͓=p����u�{�n����T݄�����B�ܜ�N�kы�wLD%g���݉�lF��|)I����t����a9��D��i ާ'�T�Iz���n'ٝ��ߑ�kl�~�N��e��i.�"i�Z�S�k?�'�etqI'���ICRm�9����θ>��m��	���CƠ�	�0&���
Q�;�A
�5i��f�>�>����ŷ9��0�B�Z'ц�^������kM�����z|��c�L�م��S8.�G���}�@z�-��
�N:�_~�4�`0�>�\{S0�H�׻�;�qqK���I�s D���v�HdZ��;@(4��x��(
���gC�u����is�0��c�yYH��1h�6�V7�@�����i�M��F.�R�:�5M���-][�Ud��	"�y�r������}�S�((M~���M�0 �O0�oO�FA�s�]�Ҧ�曯.k�"�o�Rz���c>�#��=$a�E�@\��A|����h ���s���J�@����^S��-SP���{��@�xd����X	�y1n�з�F�t!
�aLY�r�6����!Ֆ�]B��!N'0.C��bX��}�b�B�>�P%p�\B���_W��O� $jY�Έ�^-��t�#/�DA!!'�ɪ� -#�n�^�D?*gd�N�MD�G�6A�������)��)�)5K��W�Ͳ��ݧM ����"�@���S	n�P�x$��K�u����ԛ=��}sfd�e�j���Gj��ab��S�T�a���fۊ�S�9��.n�*Z±��>IY����o+.����9�uPR*�k������&i�TGk���l�Lpt��>�����7,��F.�~��ӕ�݇v쑍�����G�vLd���h%N!~�`������+�%�%�C(T!��� �L�B��g�tp�k>u�kꟻ��$�X���ҘO�A!Y�h'���%�Ϧ�b��ʞ�]i���l���5�?4�]�ѐ'k]���~1I3���7>S�Ă{���lx�)��ާ�F6B�m���3�;�40,��B�lp�W����$}�(�ɔģ����(N�ѐ��@��v!t�4�_Kh��~�E�n�?���p��8�`�27-��)�-	ۗ4�^�y��H��k�Ig�a��{�]kb�B���\?_��^ޭ �;�����m�O�:nڜ���.0�@�;��)�g�/g��π��
0�>��nR�+��ж9E�ҧ^���t�|)�)&D�p<%ӧ�9Af�,�g���K�[���ס��-R���86-.!�Z5X޵���Roɞט��s��{w�T��5�guŵ}��e��7�.|���a���ਭ�w�F`!�B<X�Տ#�M������BS���#�cb�Sv��i��R&��_�ɕ~��Lݶ��Uʶ��&X8��M���W�s�����;#Ɛ_K��a�bDC�+r�]	��r�+�Ԛ|����j6=dfT���2�ct���;�D�fp�A���H���æ1�H@[5v��ì1��:��%�=�f�3���j�u5�/V'�Ŏ��n#�7��U�V���6���o�������-j�xC��6\���iDf��3���ySCH$�ǂ�WB�����d�CF��$K��:� �s0�E���Q!�E/�Ho�x�P`�4�c~/��Un6���ԉqG��3�
�1Z�?Up0�j�<9����ŗ���G������өD�üic�� ����9U�#�z�R�A����������(�+�D����G��#�#�C��"!�'��3,���na1�$����*؀?�����7�D����l�6In̟i��c�_�G��cw�᣿B�M�e[�Oe�����?@�����7����L�\\�#�^�э,!�d�Hથiԣ�o��׫�Ӧ``�5��L<e�F��I�2je¹&�� FB��E'������IeL��K�E��CD@����\�Cm�ᛖ�]$��������	]֝EANE�
q��V���=��4�6�������m���������%�j����~S�+�⏢aN (���r�y'=��Q���yD��' �kx�����˞��Ǧyc9����B����N�m��1�<eLq�jg䓍�[\^7v^5T��q��d괯�ļ�!�,�z���	o�C�7˿�����G����6O��r�v��y�+3��� �=��]O��x����S*|�A ��֨xD����ԙC�Ҟ��PȎ/hN��
BX@�G����U��]N�>���=���(�lPV�f�S^0å�/�֒�7,��� .���A�1ĺ��%���߫ӰpM�}�ȘQ�"�� Fh5��Kp�� i3Trq�n��=0���&Q��nM��~� �=(<���>��nW��"�Brk<��4�?�%+Gʭ$�%F=U�	���+�/
R�����nM^+cQ��R$,,��������?�-�Z��<D�JF�c�H�2&�����l|��fY�9����O6[T�e��� y9������B���2�z?l���a���H�`P���UŠz9w��oqG%���%�F���: e��E�d�
��N������n{�eI�{����٬��=פr���G{�ɛ�}����d	NS2�8���d*�v@��� 0�F����}1��Z32�ZN��������B	��؃>��p�o9�Ξo�#s���/QϘ�P��4y���B���7@䨍��-7��PV�)�\�]`�g�gv�nz������':#u&`;���+�{)�;�?p���9��v��>��`s����� ���2�mW��Gk�%("%޺p'��3�ݶCN_��s>�m͌��y�qӒ��13�؀��N7�
=a (�����ōX%5��/�iy��U�G�MϜ*���>���3�Gʻ�i�Q����nAˡ��|aW{
�k�����6�s;���\�����p�p���z�䎂Z�KZ�,��u��^��h�l��.�j6R&�q�r7�*-��+8�w�9&�<_+�7%p�gӠv����+g-;�ΠxoW� ��>�k	�=	'�i-��I�޵�B񴃂�>���h��!�~㢮�ڦ�#�W��`�o��Y��cx�K�s�̑�b�\7.{0O2�+�4d����0�n�~�h���d��tࠁ�~�	�[��Q��q�N�j;����QkX�$��ߤ�?�R^	lӞ�?���Ty��Q+ޣ����/�B�u��l�<A
F�BvmP�� 0���.跇u}�F����VM�