XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���핁��';�q�Z��L3��e2������w�ت	]�ڦq��
s��K2�F�0����]{߂6����P�i�G�B���A���SM�� /8-�<H#�c�O�ʬ��>���m�y���y��>d])��߭M�E��ai�������Q�#�R������
�G�+f�M��r#N���ȩ������~ N}���R?s�ySo���[�4��)KI*���ʺM3e�Uq
�2�L�o�8J������!�L*�B~�q�o������dK�c����P�(M0T=\O6j���0����ȇ�&�m��kV'��HYj�ћa��&$��������H#c�����fC$�;Z����X!�	$e��T�����:����(r2H7����� �mg+�jQ=�m�b��o��8?)I���Y���A�Upç���V��e
�n%*�n�4r�B�HBV冚�R:{ְXn���o\�`|ٽ�����X((bLW�G�b����[��R�Nv��8\��B��yi|���MC_l[K��ݯ��bm�z%�%��1�E�N}�x�OLɒ����9��9<�!�	;7�Q%s��c.�7@^�;ap��k�F����(�p���Ǜ�;Zx�	㿀��,�R'���n!����Ǽ����Р4�#�� �x��j5�
�U�No�j �͏X�6��`�"��NZx���;�5iX�Gi��LR���F|�3��7!X���ܣ�K��!���WQ�Yb��A����SGXlxVHYEB    1853     810u�K�!������B(�#P�W>�O�M%��D��f�]LWD���;�C�k�)����f&}�v�!��F����NRX�+��\�C��t@&��,�tM�:w2W0[5�R��!��m��4���&Z����_�ؚvi�L��l%�F_TU����,0�����3m\W�. � �.�j�� �	�R�ӓ��� �1�*%�r^�K�YZ���v�5W�k�:�{�x��]��d���@��Gf����+aœ��1�jq3��/����M�߶�A~F�6�U�"��'(3��I��#otu�L����.L*o�s�q�Q�8R�>�I<@)Xv���g�9��-�R1�{s8m��n�p�D��1y�d6����nZkg�Tȳ>q�|�XQ���2m������ɑG�oWr%��P�M���k�SI�A�*�}K������RժĢ�-/|X,��Tq���^N�#��4A�O�Nc�j|�qԺ� ��B���?�6NW�b/r�s��D���E�5?�I�f��C^��Ơ����%�g�]���8���\Vm��|�
& ���*�R+�y��&�j�%�P��X����  �̷"~��3���X>����O3nۜ�vծ�Wla��T�5���c�/,�a���`�wm������F͵͌��<��bm���J���5��w�M��>)=����B�,+���κP� Ƚ0�.;��9Kl<��l�ԅ�:�0м�����F[�V�r�3�Fy�N@�;���P���B]1�͡H�0�Y�Cz�e}��0H0*�*NN� $b��X�W�q�k�s&mj=�9%�-wlB
�m��� �!t���E[�(��7���Y�U�lM� �1wR�CR�!��@� �=�xӏ;!�{0�=3�S:*?8���"�ЩF���}8D0�	qMeuoQ��U��pi�G[d����v��Ydc;�*��ct�
&�FI��=���:�ӗ��ոO���Z1y�&|�sƪ��!iB����+���\�[��S�-���`>��K�}$2O�1s9g�P-�w�}hz�W����_�6x��Q%927��%l�8m�4*���c�\r�,P �R�kÌ��W>[F�M_�gn�_�&�ٰAt[�'����lxOA2Uh����	\�P��(���/ ���#�z������uS!�l=�[c�g�Ѭ��S���Q9���U��̩'�&L�Ɠjc��-��6����q�e�9uDO8�y+�U�6��c�v^pت����Śڨ�JX Jf׬-Q���B!��4��2�3���b#��������`~O�
_U3i���~�� �կ���u�'�:x]�_��q�?جtט'z��I��_��ũίR��p��Ģf�wG6
C`qշ&Â��YǄ�yl�`Zz�M4|��Nl�� �h����5�5�zg���8pWg���gp!��7PDY����k�U�ٵ����T��5[�R3*�����v����W֏O�ޞ�/h����f��6��Hj�m��KҾ3hro�jP
Cb,�K�#1�Y��&�t呾Q�`��� C��C�j����(v�z�K�̼p��?��{��H'�)nR�g���J�g)t��pd�R�>���E]y�����e�ʊw�gv_4�J��[7T,���d(R�.�O�y� ���"=���i��]c���J����y~�z��v4���9��q����L.�F����E�Q(ʏ��T�zZi�@��u��l����$�	{�}���1A�LD.C���FϮ+�U����_���n�Us�Y��g�m���$��ҭe�"AOg{t�Ͻ��f���De��fJ�5K�^&*8[�
�Ԁ��^��0����r\���s�j����j*n�H�/�r�:�"�h����w��E>I�☆�[#$0~U~��rK#Km��;�LU�ׅ��+:�N������]U��G=+����L>����S�X��T���@�Ȗ��� ��(T��P��A^�|���q� �G{� �����9�c����Uʜ�v0�M��