XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m|:5H���܈]���j���A���w�-5H��P���؆�} �f��Дq
�!���Ş�_���Ɔݭ��H��;���|	���a����H��!i���'$!8�گ�	`6�T^zTRIM��K�L�d]'_(�������F���)`��\��G��t};s����`>c�G��[a��8�1q<@V�ն�UgE��Zb.m͝��p��X4�89�k�:h�zk	��Y)�A�ƨ=t������:�VK�K���r.�8��1="vZK���Ɩ���[j[��(n7�{��O��R8�VT,��K蟂uj�3�c��	�k��ߴ��M�a�����FōT)y��M�p��N���^�v�ds��'�	�b=��>�S}a_�|�	��^��$@��}l�V[V`��=���8$�x0Җ�^�=��U|��#�ᇵ`2E	�������흪F'�c���ݩS۩yT����V�j�G�NS٬+�d�����t��g� ]�@CD�H�x�T��SF럨��'K���Ov\Ȭ �$:��OL�ԛ�.R�yԂ��ߛ5uO���Б7�Z�) .�Ss�ͯ|�}_�\��U��b(�|��ѡ��x���0��.��I�bإ����Q8�\6��a�N���=��/��Q�O����ío	\��|ֲ�	�&��>&�ٛ�-_4�ܭ����1ɒ���4�M0�ZB��Z&;Ln��,�m(U[��q�[�B�fNlS���奭��4�ڲ R7��=�QJ���XlxVHYEB    fa00    2040�;/:][H�F���05�Xh-]G+�LE�o�%w����{YU%W��X<m�l��[y��}��;�fs�)m���u���f��*������Y��D$�ڽ�����v���u�,we�F"�zu7�T�i����4�7`H_5o��(��x�[��?�Yh�V�Y�vԩ0��L~��9�0�{̅���t�*�J {�����=fZ��g)w�Z�1���(�Y��@ܧ\#���f�vk��ˠ�t'8+r��NЀ��T��y��n)�&�J�>�k��s��7�D���ۀ�}ջ�ɉ7�!Q�4��������{�>Y�j|Bǅ♌�Y�����`��]y&Ѩ+�0ADH<�ja��D��Q��$��H\#��z����鄐<��+� ��9
N �J$a{�gn�����w87$#�{Ma��wη�/���a��0�S��ge{JFA_&��~ܰ��f-����>h�x�ݠ�g|�.�E{�s��y���	f���x���#4������6�.��"��W�Ǽ��0�	"a֘�u����ZNѲ�e�6���!|������4��aWY�+>?_7������r*>6H��̢��IM�/�x���@&�a������r�Z�����RRAT,�;�,W�N~������՛��"5x#j1rO���B�*�2Ǖ����&�O[W��}\�Z>�
�Z�V:m=����l�*�*�S�����]7+��;^tm���)������������B�񠎒FDrb�����ك|��l�!mr��s��}��0���wK�l.��bw��V:���s�\�*ADH�t��y^<cc��F�3B�}J)���	�e��ݼ��#j�=��*X��%�/�&�����o�-�$'(^U�F�S;V`qe�O��u�R��7�A|h;���K'Z������8mhq�B	>s��\{\.fElO��#��)w�\��$�Q�`��Ɏ;�	�[���_[��	�������"��[xlk�S�qv���@u�M����oy鶚�&CHy_֤t=�fΖy�O�v%В�ù�,���&� [�`#Z�= �|9Y�鉊v�/�|�ׁ��֯�*{h���{��o�c�%�.n��H�X�x��q���J����Ņq-�y���W&�xi�y:�Q���os���k�'a���'�~�ԕ�,����:gҐ����[�R�R'�'�|���D��]?�o ��a��A(K=�f�<@ۜ��钕ۢ��J��8렂�_�k�W�kg-@d�flv�Cd�ec�X���W���6ORȣ�ڶk�������!j!D@
��|���;�
�U�e��S2Z��qV��d3w�X�M�0~a0��)Q|\����n� �A�3q�+͊:/��%�%����Q�:@�-�UC<[D3��k�o�����ا)�8����'1�os9j��L�{�]�	�~RK!�����Ġ׽�4) �.�WHh6vd�r	���~�kgʽQW�wv+�D��@� l�.��O}<+��j?�<�Xs���S���$&��Lly�����6&� &�9�?�[w�����^��sr����������{�$`�T��|�����f_�\%��2�<}���.f�%�r�O$K�+����?}�r�JP�8p�H��ghM	z��!��vhF����*+���&�'=�j���u���|���;�u%s�q�'��H�+��T�x�H]���	iS]�0�_{���DeJh;��]JXxO
J�K��ZP��p|%T�<y2# p�������D,pUa;(��=	B-B��*#����$�X�j�-dǎ$����d�80�|��G-I�ou���8���8tq�s�E�`��v�y�@.�H���3���K����B?jA=�$� ��s���:�F��m�����{&D�^{ ]�V��2��Q37�h<*��]���B�Uz�����W�|W�����tja�����$���� ���p����a�gؿf.�j��*p�<���9�	������`��v�'j����w[-h��{һAc=�d����]h'���<�D����:�����'=��R vc�*�Ф���	�A��+����hп۟Z��4\F���a~]Q�3vD+����t�>���̅�)����`Kq���_�Ί��8�.<ӈ��c�43���M���He���`�#2v���p7�
5-�V5��R�s�>�a����n��;�7����{ٛ�WK��<V�������j=:��.���|�TP�G{�x��d�/n��f��=f�ٓ��6�2����?H����ބ�V�L����X�f��(v�-�}�E�I:V�{�(� ��5��wR���[�"�d���_*XDbL��/����aD2�k[%R�44U�Q�j%P<�0�%�"���V",��^3k�BEx̺n2T>�@�S/	�c��2v�W[
�}٤=��[�[���Gq�Z��3N�yȣ������V�Fz<æ�r�1���oj0n�IќI�ԗ�ط�������m3���`�Y*9���;5�Z_(k���y�a���竺��4�s�K����0Sp��7��k�<��5�I�[��3Ĩh�Bc�D�U���j��a��.т��|�����!�ER���v˲��n3�LM&�"�J%:::��j.CWY����'G���YI)�`��6㤠�MJdy���%Nq��9f7�0I���i@7��t���A����J����O�5o�W��FJ]U�9��yU*�|N�]��^eڏOu�Q:������4Σ�Dh
z�8�؟��A���������R����6D�q��q#	Q嘩[w0D��FH��T������n��\�7<�����^{�Å�~��О��y��\!��5pt&ȹ��(��hg���:�*�{#�W�������ھZ�Ss���㺓pf�b}�`ύ��`�ꁔ��:��H���E�ƂV��|��=�W�oF�[�k������7�Sye�Us`���ӻ�!��H�����}J=�<�c)��-	�5&�X*$G&8�:'�m��` 5� =�eg�f�R�c�X�=̉�{mg��>4��Ò�,�ecY�IDAD~��石�ב�E���1��v``cs*l@�u	(��M�P?'M_F��ښ�&W��]0t�!��� �0�V�!�^��a��Ѵ��;n{d>��p�ii�?v��Ɉ��_*�{s:��c�H���uq�)��� |�5����Wo�9��[}�6'�j�kg�;����Ze�8��Ls¸�ݻ�ry􍫄�m9���O��� rS�Rg�{"�K+n���)�}�"��w�b"BXk���S���l�k���>��cg���j_���^�4]��:ǊA�ҽޏ5M���ڋk�!�Æ���5	*��U�����w�����S���U�� �׼��	��`D6��Px�H%�������S����~��!(!�@P�)��⦪�K��E6V�H��5P��bMo�i�a�r�Cs-c���O�M����!U�/���F�!}=f�`y}傊�!��i��i�g�iŇ���E�w/��۽M�\�,�Z��:�1V���f����ȍ�O�1ɨsՎ�B�f�(��6�m �z�8�R��е���+��QY֐�]4\	��$1��<���k�,�a2n�X���_�E_mMSh���w��5~2���VU��ٯXS�Qg��Ư�2�*�LV��#ݻ�Op�fbU֠����ֆ�F�~5�Ϩ�����$$�H��-Q�;����o������$6c@�8�a�DH}#a���9W��SpR'��D�gK8�N_��\�C�QO%�K�@�ք �Gk	�`�}�n�;I�^��7��.ѿa�ɒ
�������p���${{>Χ��xfS	� �"�p撩D/�Y�
Ƚ�X�wF&h�S��a37��.���,������x�GZ/�U`�n�X!T��()"ɽ��zOÖ�h3�,H�i!Ӗ�w��+,���o`R8�^�_��x����i�fO}>!{�N�X	�U��7�������.���r
�����,�?�l��"��~=0s�������R �p?���v(쫸~��[S	95���
0����U����DW \��0f���%OT�u-�אo{�L��M��#G�~U'&bs��[6��D	��J���+	��g�T�+���J���27{���I	~j�c��u@� ��W�zW���IV�^+k�=:�d�g��qV�:͍��c�*��/L�=WWh]D����r-��,��8?ߜ�$�j�@g�QB�S,�o��|o-�JC�dx�f��}��=h��m�/G��'W��07�u�K�0���/PyPJBL�o�͑W�j
��v�齴�=�^���#��/ �J���qSy���}�"��EIN-�=ra6^��.U���v6,e��/h�dҒ��}~^"���}أ>��֝e����YٳBO#���fc��wǤ��t�����-�����|T��
V�i������=���w�ɨh��Sg�t���{�-��P��BN@��z�V<�o����?�� i�¬����|���bbz���!y�j�~35g�k���O����F�D�Ug�X���f�g&(�Θ�	�p�#�2�c�\/�����^�.=���#�Z=��� �|����/f>��f���5��3�E�x��6��;Z��q�A�"�����+7�1�N$Ac f�cF�ӝ߇���Q�d��� ���5'�����Eo:%��`0�_����e�	h|��Q��fX�6$[�e�j�ߝNk�@�'@/��K��?(J��lO�w]����a��D\�8���6��."��# �P���޺d���.�$u��"���L鬻�_�{铥��:Ճ�:3�-�r��W+ԝ�q>��v:��kmX�j�^�[�c���t������  �\�J/�A�B- ��vV\���u�fQs�i3�I���7�͓C���R�}U�%Eٔި�<���ܡ�,n�"�9x�ʢ~N��%t�1�А8�����Wl8�9�\X:�8ź�p�r`�
�n��πr�%9���N~W����@L�95ֵ:��q藍c�ϭd�����{���C�S)"׮,27p,#���*7��:a��F�z��5�]eo;�����Ib]�S�/ T�v��|��!,�W��;`���F�/?p���V�#3�5 ��]��C�D�&��8ۡ������ٺC��AJ�@6�E�Q��+�T�3��~p��Ew��x�d6bJ�	˦�4P�1�t�2���d;]�T�����,��+X�=\I���h��j�4t	b�r�k.����V�=�1�'�:��".�/E�P��[�����J����f~`=�c��mɩ��[Ty�Wy�Q����
��5�jހ ���*/ꎖ���vOH#�V2x( ��c�JG�EO�<7�SY��b� ��sN��y�5�;'�4~^�4�摀�{f�4�4NI��J>%�/-��"�")��E�>WP��f�:[Ÿף�LL���?������c�tt����3*ش��R��Y���-�8�c����c<o_�.H�-U���I�����I�b�xP��ŇRʓ`#��N�[7���[�Oo_Zun|[B��Ԩy��=�xXS�02+.�Q6F�)�L[�}��A@�,������}�9�xN�ҿ�W�ZI�MM����\�%HM���Lv�����(��R�5�pӴ*̐�U�G��,��аh�n����6?�4��V��ܬ����G~+��|�%�UEn��M��xb�0���>��ΜA�k`m���������&q�TEs�mؠ��BY�[b���κ�3O\�;�0�N}�yʈ��	׻��9b3�+�m�XAw�N��j�Y3�^t�=qEɘ�a_�nߢ�Mr�z�#w+��c=|��L�CQ�4 ���YB��\=��|�o���MM��P@Ӽ���a�9��{1��9��/w%EP�Xy� �E��K|��+ɛY�U��d~e�hc��<kD���F��@MmGX��Y�w
~z?�a�eo	�g�B�s���{�mH[J\�ϣ1����B�����=L�����@����o���OV��Ğ�+Y/o��ׄ�3�{��������W���:��7Pc���h@�)5��8]��iY�QwNS�b�%�W5��	w;ؒ4�C������/�/MDe�J+?cnB�a��@����> za��ʃ~��y�� U:�J���(�z�ƣ(Nm�}�ќs^����WEp{8����؏���wO	Sş�ef�n����8�:t���x4XJY��o��(&������}˗�m�X���%C#��֘�:�̗�*�r����=^<���f�Q{!'��TS�$�HP'sz��n�RՔ�ŕ{�GO	���u�����q����jڭX�,�������É{q?����w��Q�����t��$<��=ȯ�Ƭ-�g�`��8�w,Z-��>�C#��I��Jh>�̢�����G��a�Ժ���N[� �O�hĚÇ��1��G�E #� ����X�ը�~9�T����ڎ �e_\L��AmGg�KP�B�H��z�Q�$\��;�D�����|W`@؀�hyj r�byKB�*"=q��\��+H�At4j������.�U�z�g���>������G|O!�}t����b��f3v1��� G���PKa��=�O%��_G��o�U���z��_��<�׆�y�����ׁNQ5�����mF�����$2�&¢����8S 3�F��[�z��yV�YW�N�r�>hU�0LG�!+�MX}�$O�wy�//�fJ�a+M�m�"�-lٳ�����
C}�V��/4�IC�<��|G���Q����r�HYe���E��6�p�����F�p	���@+��d�m�H.HcnZ()w�,;���qx��[��Aԃ?�_��1�Y�g�bT���l����E�F�'`���;��%�-�^�?��P�P��o5�����/Ϩy��7ڀ�2��y�D�Z��	z�s{�����@�hy��m%�M����w0��^;�ܚ��^a�Am��T�7���lPG�+](��m�D`TM��-Jbf�P�ߘ�w�� �!�}�$E��N���~Y�Ȅ�c�Ű��Pum���Z	rbey)��+��ȰpS��24����2:�o�J�?�����;aD�S��W����.�!��ϳ��AK��`�@϶�);�
m�t�]
z����T��ׅ$�X_^h)m�?��Жj�U.��7fR��x~�Ķ��B_�9��D��^�TYz��$@K�5�f<����g-dW�e"B�Nv��-���[��C� �e�*۽��
�ꆤ�)c2�e/����.�`�m���}
�}�*ڹ3*[��0z�q�%���O̥P�ta�X9�'��|���u�*5�Nũ��9�Dl��8�+*
�A�/��y�"�֦�L���V��kݞ�na����Ð?�&��Mq��|$�<j�;>?d7d^"�p0�xi/?�(�A���I��p���Ly4��
7f�P2 / ޿IR��"��ٍ�x��~s�H�1���� �&q]Œ�D��॑�a37V�t�krύ���EJ����f4ĺ�����'><�9�V�)����~��(�L�hDG�b��	�90+-�X���*�d������]}\X�"��M���e�j�X���!�$ˠ�{1^%SM�t���␸�6a�F�n+X�����,�b�-�j�	a��C �A9��]��(��sh����B1KMZ�^�'��wb��s�V%�4�<��T�DY��g�Ǐ��~��^������y|2#�|�$���gZ�PC=�D�r�K։7�>s��-d֋ �'~v�/��Ѷ&���i ��4O��%G�v���XXn0	�u�D̎�յ�?���I��C���(x6��t��R��*+�<���պ���*b��9���D��$t�9�L��wJ��?��(����y�i��鵱5�'��Hx��?�Yv��4K��uN'�XlxVHYEB    4f62     b50����,\��dn�C�n����T��㾄��ªy-��ܰ-�3l��'D:��*[���mz�;�-�??4��-��^�<�~�[�W�c�t�
�|{}][}����ʮ��J�^F`���j�:�(�O��<����I�[u~��/d.	G*�kmBzL�df���x�W�s,�ڳ� n�9��O���g�o�[�i�{��]�fASA��q�4��`hQ��U���b�)���l�	���:�0R�Y�;�[a"�#���=i8o��Ǝ�1p;ݙ�)Ȭl"I��է�4Ƒ=�DB��BB
,-f5�,�Ai��=*>��(l���+g�#�P�
�:`m���ӖLR8x�	)�␐au������Z�X[&��d9������ȑ��<eA�I_���,�df(�Є�i�¬Cb�F��i�o�R]K�ć���N��lD,�)�n���MOIu5rORɸ��0�o��k5�<W�V$���>�s���ѧ�j�d!k>��#%&�,��KY�uG<��\�@K�.�+AИ�ǵ��	���D�2�R�zB�o�l����3��=B�?�A���GS3�d�4�< (ؾ�oS_oý���~��@�ȉ
�/��XN0ife�#�-�[�T������l�G��Jr�m�WIB����ҁ���H�-(+�<��e��f�f��?H����\���o"��=�\P�����۶��h�B��Н�֏c�ۃ���/�6΢.�.@������	z!����+3�tΝh#�aC�����E�[�8�Nڊ���?�ǁ�)5���d^��>�Vˢ�rB�C�@��4�o;��T޸h�̯a�#l���&���Fa��T����bN݀�țh���mF����d���
����0j �r8�ҌD����8=P�
<�v+߳���K�ʄ����OX^R���mTB�tL��R��ql���`j�f�8��.����QBzvf��������?�PZޒ��
r�>m�`����Y�N=�:�>�Cj�%z� �����Vc&ɍNN�a`���Pc�N�b�sz�H-N�ZB�h���`�ĝ�H�?Q^P9���<u�g\x��jfu���a�O,z$dӒ� D���\@kH��$x͠v-��ډ�q��j9��~L�	D�3�iY*�)7��D^J�??"i�ĸqu��3��7t,�	��o�q��<�Tծ��Z�t�y+7r�iש�!�X��x�H��(�-�ޛ��߃c.�#�}�5������ZYQ��W&MkM��,�H�D����?Ȧ#q�B�\��Z�����T"�.9�h�#Hgi��.=�^����c�N�f;���>y�J�$>Xr^�cX�L$���Oo�bS�S���|_N^���� ڤ�v{��9�Q�l��e� �YI�u�09�Œ͆�Ύڛ�v(�>ߧnN&	�M�a����A� �2���(�����'=�Z{ �]�،U
|Y�r��&�!��H��ݼc����q�E�	ھ5l�4O��6�%���B�Z�M�y��/Gi��]4�XO$�)���{���v}x���p�ӂ?�SH5%��훚 ���E��G��J�-�\�4b��t��ѺM���=e"$�ݧrJnG�X ���kc���9�L�E�z'����i���g��S?���!�,7>(n�:�S�̀ҍ-�`' ���DiG�{�������Ҭ��ܚ.:-R���6��,�1�&e�<�,�,S�.�@lO�uT����oU�ҫ,�D����/��t����TY���;���Bl��S���Ƒ�f��~��N��O��OW��Uxy�`hg���)I����5~���Jx�y�;�,����,rV��J~����?������̠��rj�עވ&;�E\|!��W�P�>��:+����ZUQ��9�L����f��}���gT�Zs��tH7%
B�ݍ����#��K��p,��<I؍��C\�#d�KW>��WW5��:�s�>i��7�a�������3K3�3T�oba&�׀�d87�mߪ1j�]�i�m�o�;�H]UDI\Y� �S�����3%fu�Z�v,�!<}kOW����s
 cE���:�ƫ�*�g����g+S �ނńՋ��0��xg`���O�]7�x�GnAg�){��anl�����ϣ��L�����z��Ϸ�5;��p��/h�6��kj�*M͵Ev�34�	��R�
}�yރR�����%I���l�c* .<[�}J�\�v;�����?j��A>ٝw4���;򢇨�W���"E ��?� �&�q����ٕ�d�;�+7���s8��H"W�#8�ܱTR���J�����թ���[k����Ү��ւ}q]��#8���.�<dꪮG�Ge�͕��dgF��^=ĩ�X�r�k��Va|��/!=�)#�Vh�K���d��kN�2��^�]�V�w?T���[�
�>g��9�A/(�r�w�*�;SJ���eq�QY+в+�Ut�/ER�nW�t~��o��H�N�@`���h�X�Ew:U4�b�ߍ���f�i8�6f��[H ��@��G��Ž�"�g{�g��,��81>�(�3�DN�m�+�Q���םy�3�g�ܷ�b�m�9a��v,67�\�<GD�UF�������hL���b�#����X-Y˷��N�5sr���Y[��sR8Eg)~͕3#�fs=,���+�D��xD��Z5�Aɜ��TC��h��R�@1�b:Upʏ�g)�����9ږ��a����+��L�cB�i��~�)EmC���P��W=��f*��Ÿ�H�?�������if�c���ٛ}���c�m6?u