XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B��`�o#�S�TQ��SzL���o8[ n5��Ml]��$;��,��Tf���Z�:�"�^G��V���4�b=��WB���8�@_���B�	�	�Z� ��QD�6�(�i��c����U�N<Ʋ�&���]V�:�~���E����0
g��)g|�"�l4�,Ʊ˧z�U+�F`�C�:+�����*�d���[��|��|�]#��<���X��d	�������o�@`y����7��Y�-�Ґ��S�5v���	�{�z��(r����<�����x���H�Y(d��˼�ZN��٦ȁ>.`��X�Z=iV��T�%��VN����]g9�V��;CdZ����s��4?7��7�&��J��(��ə������Z��RG8ח��.ʿ.8��F�j�l���al�Mj��:���p�����eO�խ���3
��=��J-*p��8q�<(��ǉ��(0�8�ќ9d}�����O�~rY%WQ���H���>��2_�,�q���̄�=\E����){��©E+Bx�x�~)�0˨.�lX�r�m������
:Iuw-Hr0L�*2�]�=�|k+>��u��x "l2~��wE�).��o[c4�](�le7�K���ޥ=�+)�N��W�\p�$�l
{�7=e�\�3iK'��G�a�R��#�{x����wP2ۭ�1j��W�M���$���WV��;����1|�2��.!

rV<�Ғ�lD���^6p�|!�A�<XlxVHYEB    a037    1fe0s8����G���N�Ҏ�L-��~j�؜���Q���'׃Ny����j�v���o�,�7�9W�rЙ�7-�ݦb���A�z��ڛeQU����TOW��j��Q2�J�tD�s�U�}�����~>
���<}���Gր�&�f�T�0e�#��d�2�<�2�l��L�M�Z�Oՙ��-F���5 �WU�-߼��u�^@G��/�Y��
����#���]�)�4n&Q�C�:���]�.C��m�]8�HW�� ��?q�����M t�H_K2-����L6<Ը8Lj�hh����`	Mc�o ��x��R"�"�� � �ڂ� ���T��C?׼�7�j�A��h�#�ڨ�ES:���!!���� ~V�)��^>�[���ۗ�IVb�r^����j��R�L�zv���[��h\���5��z�P,;�Css6�8��Ъ�}h��W�"~��-�
ͪ$�6�a���i�z�-'��,��W�^i$ĳ��8c��Vo��.;j6�W5�����ڥ�Q�2(�E��U��^S;m�nz�4�W�˯0��9n��o�Ƀ(����خ��o������r��#
�N=�O<�g����h�b(rM)>U,�;����P����?h�b~Y��,�G.E��?�a�Fg��rd;7|.�W���8�fe�9d�1�:�d��]Bo�\$]�j"�DΙ*]�/f���;�Pܟ$3���Jr��|!#g��F�EJ�d�ȼF�D���sڹ��nN��>���jOH�±~������+:��"�4�[������E*�Q�eۥ'�&�����?U�v�%ڔ/� G��qE���66��~����� :+��W�.�Fޜ�%C"��W��t�˅h�&���ԯQl����%')�:�o����2鿑�`���P��g��A؝��F�6 �|_�>k%�"�n*;��A�P��і'���Tx�~i&�<wȫ/0���h�z�#��$��S�|�`ѰP�bt��MR���0�@D1���$��9�nln[Q���G�Ȃ�)vzsi�Ч�$����e#���E��$��(pU�s��qV�#h��}DD ��>g��hϷ d���I��Vlb4�)Y������'76DGM�\��������:΋�-0L�f�!��<����%m��³ՠ
�y�=��u{4z��N�4�+���G�ݏH�&���;%�g��j�G�qb5s��F.@\����������u��;6��Љ�{�(��wX�c�	��#��j����X�~���{1�{|֦�h���v
�[������Q�1&�铦�H�HV���b��QC��j'�$�6=����8 F��3�n�V��ztrc����	�u�c��V��_B�� e�Zv�&F�?��Ў(�2���+(Wօ, �t��Vrn�A�g�||�uMCM�J¡���LR?7�)�b1k
��j?'Iܐ��.i�"����Y ת�@��˨������3H�Ƿ*/dC� 3D'Yg�t�#��FD����]��ui�돴�Q�+�w����N"S�ڃ����DF�&U��|�N=���|��I��m��s�V�aڑ&$�%P�S�����ܔ��,]���8�y��y��6���d�M>��$�0%����������
0� <қt"��5�L��T��T��6[3��	���<31spa'��;�.Ū�0�}��I�50F\Td�em_��-BB�#��K�����?�`���	ٜu�����ٖ$bW�"�%�Ũ�s��KE;�§}f��x7���p���J�Ҥ�#����E����?����I{B٘d��C���v�L��j�"�[P��V�s��O����b�Q�⬶�{��nڂ�lG�_��&b8) �9F�i�����5���p����-�:� ��D�-�����G��1�cߗq�)7�O�����h>ǵ�R���n���K�L��_^JD�R�;K&��#
Y!F��q,�=F����Y�ŏ��!���6W˪�t嚬�4|t����Q�؝^������^$7S���]3��U��B���O$�Vo���h;�{�[*BKL����q��f�<0m��/-�=D�Ǎ���z�uU�T���p	x!H%��n��N{���]A[5�Q�|�z�����I��-D�Ҁ��B �;j��D��m��+�"pQ�F4��(�Z����G�����	�E�t���)����i��"��ý��l�:��&���8
��$m.{�������!�:�4�k���Z��hhU��de�7T+퇯2�~^r���l�:H�N;�F��v����M���w��Fɳ�Ǯ8c��wF�^�ˡ��t�sai�p'�O��|�AVF�
�	+�9tA���VT�j�$�ϼ�xf����2��T�O\����6���N!G����ݒ���p
�Ws�j�ٰ4$��*����J��O��d�̥��-v�l�/xo���	p�ә��^�����Y|g�'#��2O:(�ڠS�_M�DH�sj7~�V;�_���f�힮P�)���|�Yi�ʎW[�/_��G_�|�T�4`���n0�M�!�G�����Q�Q�XE���d\��S_�N��{�L�ըM�0|�z��]|���p�a�!�$�#��f]��W��
�	\m�:� �V#�ׂ�G�����; �}ƻ����	��{��c�(�����c����$5!_�ן[w"7ޱqb��ƛ[��^�5]�]e�o"D�{��2wL�An�A0s��"�ժD��K$�A�F�1�#'�YZRG�l��%���a�ʩlj~���!��Z�_dX@�ˮY_c�O��L#�t�F\ym��]9�i���?u�J�9�[�l5lHFFۀc�����0��K1�x�7�N�+��z޿��͔
$�%��%�u�? ޔɜ�~��RiYz���ZJ�#�6N(���&N²�[��
I��C��P1~Vĕ��w���8�ND�$����>r��v����aO;��!*O��&�e�dr�� ���C�c����	��w�1�D�l�~{�*d��璈�oE�J�w<���r�[��4�[]��Us����T}؀��ܽ�1qh |��۰2����+HG��"Q��m�H̚}�Wê��`Om3U���h�7o��g4�L�=�.�6��}�l<rz5(k�rx,�%��&rr�ܳ! :Xb����?���K���u�F5����Q��"�:q�R�w�n'B"7خ��"�4cq�� ۠ag�J4)/8�<�Du2&�UW�A(��Nv�!�s�> �}�a����^���V���a9k�@��o�r1E�?jD#�������c��xAT��Ki��e�6zĩ8\�~����1�~��Sڗ�eb�� its~��N�~u�wS�C���ߨ�\��p�4�[��&��E k�����j���7�aƣ"P�5N#
d2ehߎ�Z�AN�a{��~�<��A����s$��Ҙ��4��	%)8%�V������b���VM\Ҡޙ+VT�tkh3��h��'n0��7�L' R��w(F���c`�Tw�!�CD���F���KX6p�G�9�m?7��`�K�HL6��r����Xm�9$��P
:W��i�簔�n��>s@���4��U;9��)N�����Y߈?�##�n�1+�n���pLh���!��
OY;ղ�9gG&x� Nx|��M�C�s��p]lY�G�8�������-�����>�{{�&wX��+}jTɶ���E���+��u�YP����"��;soY�C&؟;�ٌ�9��	(^t��z�,��CO#��D�nQY��I��Y%�(�<�)�D�1֙Z��3�$u�ԛT����W�W�u�q\�2u���	T!�y��H #�)��F�\�ï���O1��Z�b��/Nd�^$�{߹2U�O��0Эf9��t_��AL4��;8?�K�R4����%ӹɫ���Q����G�F=~~B�>�� AN�Ā�L��?��� N5u��|,x��fu���^Z���{U�㸸�kpI��>(��
6u�+m3&�=��-�ቛTHo�����'��#16�����h%	�Jq9}�5Ra��&�[�����(/��^���p>T\�C=Q�j#V�z���U�tJp�&7i�Y�q�01.��
r�$��2�-Eq^�$�C*+��-��Ě W4lN������щy��Bn��D,�}�����t��C����+o'���48��9�J3&�x�'-��n��K��(�3 b�~R�Jq|z �7�Q ���p��w�`�1+I���tKN�ŏ�r�H��x-6U���n"���*�`�����]}ž�FzG3qю�N)����<�ú2$$^}�&�!�ǭ�'�P�ٍ,��&��	���r?��JŶLQF���������p�A�IZ:�զ�g����T���t7u�/}��әA�l�V��Ɇ��*��������ʥ'��IS�8�o� Y�+�:*�M���@��HY�{JgC���	R����B������X?�+'H�!��S,[�0zbY�r���,���4)��r\���U�"�\��-� �����+�דC���Z�}]g���%A�.��a[Rmo=�n�3
�$�8Dg�0���8�l���L��fW#�k��������:A�5����Z_��Jx9ø$F3ۦc�h��>�'�@6�7��l��R�#$�=3w�޸�H�t���l	��	���ß��י��z%�m^�.(��#� W��8���$��c=��������F�闯�n��_�]�0N/�?O��}�T �}^Ӽ!�[8��ɖ����-D�k\ٜo���@:�F/\�j�6��x޳)�����D�%lE�ZU�t^`�Z���N�,���u���U�=��[qe<NqN��lf	L�lMHG��ɇ+)hyPnZS�0���b�!W}Wn�����q������[@N���@��\h�!���(����.	��8��:�?lk8�!=�/ʭTؔ�TL�BOGA�n�,p���_ -Ս�nՋȢݘ7T�}������W��+^}�k��+z�]��jY��0)Oc,x��n�Ͱ��Rcf\��3�Nw��jN.H�	jI�_��V<V:y�`� w��=�h0TH����*�mh���ۯW){n�} ��l���8}� ����-޼�)W�]��1��''U6� bӆ橧'�.��e����Ͻv{x�7$�Z��gש�H`L-Y/��ӒKY;� {�jo���o �HЭ�/eKdK�]��g�eb,�Bc����t��~ �t�B����^�NI�ܷy����}+'k�+�dR�9䶴�ۿ7}k��r|�[<x��x�.�c͈.��BȰ%֣Gm5��K�4���Y_����C�^����5����S"?�9���/q��ap�za�.}~׺0�]5G=�zq�X�:�P�D?d$�����n��no�,�w�@b�C��Vi>0.c�i#�{W��W��蠞CN|*^�,J�'����u~�g%,�\����8��疆pb��(s��2��'���38�)*1Vk�S�bS�T�J}���-�3�Ճ'H��^���n�њq)��~�-�u�����Οp����8XVN2b�e��%�w�|���C����sy]	���� �X���T{[K���φ[��q��QᱟFY�"���3�d�Pv8�g�I(с�3����El��4'�>��G����mKKMK#8��q'C��$
�^��� |tK��i�S 	�`.fX�p���Bm+�QtY\e�����L~������oh
�K�̀�G��$ϓEw���ni̄��f5��T?_���e�@X���2��(!���ڠ����]�˷��vvk���e�H���ݧ\I����9�\���|I�7�uv��/�G��}��%�Z��7�[��8ߔ�8/��@5��x`�zn��"�������Ģ��`l��Nu?��
;����W���/��<HE]�*4D;7��QgD��e�G�Мy�`�y����;5n�.D��]|���h�X0mzP�47Hy�8��~D�R��✓����an���X�Y��p�g�rIE��Bf��a-\>O�� ��5x��4(�e "~��D�_b�$��#�r�>�=�,��y�A��,���a��4������C����p2�j��̙S�Z;��._F:��ܰ7~�y�F�06��u���j�b�e�B�eE�[6��,��(`P�0�
>�L52��]C��>���ĪQ�_'����ߨB�@�V�8���l��7��/�f�UAhz����p����6^�>�����%@쐦*WS�rŮX�P{�k�s1�1?[jR�76r�Z/�  �\Zu���Ve�i��^(��:�VX�&^[�ךr����'�k;1����ƕ[;�x|��}��\�|���l�[�@������a�y�+hU�&m�ܼ�-��_##Т<�nV���"���6�6O� ��K ���q�s��(��\�ΐ�$-�T�(h�J�_�9oF��?�L���c�'���I���u[�j� �EPe]�-X�m!,k�}�	��[U)��&�Db�M6��&�Ŕ�ۙV��`�u+]�M�����-�ŕ���P?�]ʬ`�P�V��\N|(&�y<�Hn��1 10�D"���Ԉ��ZCq�e����=X�u�$��|��k�l��6�d�ϐvq�*�dD1�[b�����=������Xf:}��EIz=~j)W�é���3C���/�g�<B�J-Gi��MW%�71
�8�*>e�q��A� p�j!���{�$��[������D��b���>�S�x�K�&���D�u��=VR��ދ��YF�N�e3�y��'ҷ��VB,��zUw�5$����8�kDåL���Ќ9��
���9��+���Ңӹ��g��V7�7�_:�j���!�)�Z�� 1��%�R���J�#z��
����~�	���}7�a�=��d����<[�oR�0��	5��e��,�.�M�Y�O�A�Ԙo�Bt=�b���d��p$&���;i�u%:{c`��q��3#o5C��%q5��l�;BΟ��������Fw�C�sh���~4���S 
]�@����[Q��� ����@տ��On�zK�:��!t�<>f�rQ�V���b13J�Ҋ��:�8��Dq�p$f������W�=����5@S�-����~ɳ��T�E��!�'�iG+���,A��V
��%,]�n�nѽ��w� �j/����Lw!MD�8Yk�����H���ܜ��D�#���W��̾�[�����]����vd���Qr�5Yѯ������2��Q����A�m�R#5���W.T��?����ns`����!KX,��������޴ZE����s��ԇ5Ʒ�l��gm�u��)��C�B�s|Fя����|C����S�0���Hw�$��D5��z��cQ�
s�y;a�{����0��-�|@�=k�}3�A-p���.��?�MmJ,�Z�(�tY���
϶\�<̠& BiX�>:8W�:��O6<;�sLU	�*.�z�e2hѼ���8��>����b^�!r�`V���w}|�Q�c�̮ט���?�������M4����]��	���)W�8��i"��g��+VG��6�@M�)���g���L�F��@�)`3%i��"��:t�<)��2��em�=u��蒸w�^��T�R@�0ѱ)�'���qcKG	6@��CW�j�,�Kc�<U�<_�8�X]�J��I~�$�o��kTet�o9����u\��q�!;T㽥�y3���z�:��1�J����%i�p�l�b�JU�Zl&'�݃�)�K�"͖��0�rH:���~`����5�^�gߢ��1�?m����Oy֬���Л	PߦH�gw:�J����D��|\