XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]���KZi�P��u]X��d��u�	�l�XQ�NGPl�,��Ґ�3!L����W�kj�4Ѽk���������x��p.���D*M�˄qd@�_/��_߈:q������P~��ɋ)��{NT����,|����#�8;��{���rF<���Q\ݶ��N�QٮZ��c*��0ru ����;T����M�YX���3Eυ�I��9-M&r[� yI�%�0E�Z�� ����+�C'�#�fNAc����ZgUM�Hb[L����j���m�d[ �8��ǦsfD�fb)
�v����%��H;�YH�Iv䡍�������]bq�)m#��4XTV��8��.a5���Dc1�r��yBI8$��Z�Ϙɸch�-�Cۚ�f������vxm,ii��Z@�(`���Nڏ�~I�<���<־m���x�G�e�����9%v=d��Е9>������ف���6�cG-ڹ�1�)��֤P5/��-�?9���K8�(U5U��'����+�꯱��&¨A�5�aF��n=�~`��,��L��˗��E5=. ��y]YL�z É��3hΪ��tu%k$���9n['0��>�����d�?�.���`��ʁ��O�D� 6O�# ���ZdK���kf�9y�.�9d;��?l|!mbA�v����5���S=. �|tI�s�q?H�����V��Ax���T���{�+r�-�;���@t�7�DHh����N/����o�Ž�����{�Ɏ�35��A,bXlxVHYEB    a037    1fe0W��~B\�Ľ絨��n����AS�)���g�c�rc��K��٦�A�g�5��%�. b�p}�?�
���9��&-4�����,-�TMPf���M�t�l�
vK��T#��s�1��4W%.�}�4h*QN��r�?���(d�85.K�h�e�G-�����	���a0��>��@y<�P��)��Xc>��[-z��n���VHx�[r�y��et'�׿B�( �����5)�=/VE�����*	E	,�I�*�S��C@9��� A�CS��6�1e��������hi�J�k�5�v�"��9�-�`Y����=ځ��]��Pk.�\6�2�A�"ʓ!Z�Q��9%�����U�
܀�E ��&�?C� FO���E�:�׬�;��ZE�����c%����P�7.0����Я���{��h�C�>1V�d=
ڭ�~�{wK�E~#窟��{|n
3݋2�$ ��օK���BD���b�5�c��\�W^M�	/�y1B��غL�Q]O��D0�i�0ĥwւ�g��͗&��[1^$>�:�����x�Y1^�s%����%ܸ6�S��c�Jm��G$y�m&^��k��B���p��OJ�6�?GA<��nH4'<���(]�U��J��� �*4�i�ߖ�E��qkp�3S����q�*(yS����8�\�B�-�IkBoo.��N�v�y�:{Yjմ�B�5�d[Ƿ�5��+b+��_�|6`?y_�C�l���8] N��3�:j)��:'!ֈF�vK�L���Zz\�Zv����c��!"o���n`K����S����G`���䈥%.�B�O~�{��[T��Ғ�7��N�=�mj"L�]t�\����^A�ܻ9R-�/}��3S�P��ħ�O�b�O����)���H�S�l��z�q�<\������q�����E_�iZ�x��kxl��<G�e�/��P�4˕j���m[�� -Đ��ƾ�NMSy�n�~��9��x ��.�a���CJ�����Fk�Z+w��"��-����줏� h��97m���3g�$
;u^V���f�Y���ڶ�X��^+M�k���rv��́`��\6�A�xOd�I���%�:abB�T.M:�"�c�#%��)[��c��J���0�h��8^޴����A"A��É߀�b��ү�{?��#��X���-[P,�lwyR��j�9Ą�&�<�� ��stf٦�r���[˖3%w_�MF�D��*^�+���[�u�\�fUW���|1k9,��g����7�����,��2�5G���^)6:��+W����`o1�CN�~*u��-�g7�[R���A_Z��W������������'og�щp��fXJ�~4D�Ywq�&VNvI�Ba�/c�loCc^�`d�3�vY�<�g;n� ^�L��qxfK������V�;`���I���J�ܲ{�?�j��(3ଏ-в���˵��e�h^Yҋ��]���'[�HE�� ��W���V���������_�ྀ�SVg�� �U�dV�T��Z���d=�,����`����hm	����Y�Ĵ.�~�����|������O�S�h�+εe(����@����7���ܸ�]�Imӫ���<�t����ӯ>;�<����A�����F)܂c�g6;j8%t��3�HY�$��«G�R��]�b-z n���<{�a����}�*�J�l*����ϱd�g%��(�j�F���9��KWO �p
�۝����0L�tE���0��ƭ��ε�F5��UX�-k5�������$'>9II����*�� �! (�����t��k�"mM�����o�?���ʝK�N���a_�Iw�&A�8�qo>���b]3�5�o��h�C��!�|�A�q4�����6�Xx?w�q�;ѫɜF�s�|'c�« fS�q&Ԟ�uFL��#	g>��J7os����*t�y�İ=QK�9�&/��-t�=�y?�F��7ś�8�[�v3xl�ƿW9�t�D>YD���N��	+j�Y$�����T�:Oz���m���]{�ɷco�����;-HW.?�i����۸+�@���	.��r-�ކ�*�2����F|��=,��/<߸'$�&׍S]�\td���3�ݿM��I#�'t�U%���#�B�n]��Jxއ��������C���������r;��Ӱ�k~v��S��ڈ���G1�ȃ�!<$A�qIޜ�֡���{�G�Yl]�L�Sd�PC���ߘ�����6Ç��B�U�rfPѝ-GU��
�Q��;����J
���.�
Rl�0D���]9��:�V�O�ÿ��1"�O��9K�2[��z /Z�46�*hO=&�ֆ�<�'"|��)�X�s�7Y�+#�Ʒ�/�K�g�w
8g���?%�Y���Nl.��;N>� Q߬n������rS��y�X/mF�NX�}��%�K��[mPJ��9ڕ
e��iY|ӥ<��ucX[^�[�̱W�f�%��pjO��}Z�?�>�"J�
%�4�I W���~�?��p�ĩ���omV���d܈�;D���������q_K^b�g�p�ن��?�a�:�N6�9�o��t��-t�R�g$�5�GS7`(�CvM�bA���+ɆI���h����`Q� �	b�i ������l·iUE�W�o�5����f��&��t>���pk�������s[6���ɹ�X��v*�4p�����?�-s�hE���{��SFq,1[�������_����m>q_���=���b�dVE��;n��1�:����]���w�\߼��1�ys�2js�y_d���tK�]��E��1��={�4Wmko�8�.�@����C�:��J�Ǉ�U�h2��/�y��������t����ii��ʭ���q�� _Ij"���r�g-��QzF����{!k&��K>X
���qLD}b����|�.{�AO��\��3P���]����޴�z�&�EE��)0B䡂���V����}\�Hs����� ����6���T?]��A�v��-5�$6J�[s���{
��>�|�S��/��f6=;f̎��������a��e#�dv+��Y*W+^��Ɋ���78��$� �E���@��H�Ir���S��j���G�;�����njwb�D����b�����Ohh<��S�Ֆ��z��
!C�jYP�A���n�y�{��  �g��9O����Ol3
֓�ٲ�w����"��_�)A�1�DA��� �"��X��Uw�y��ݖJ��������v���5�].]v���.c���\gyk�|�J2-;�2���"�ٛ[)�mA!)����Z�DI��f�XP'�#��%���%>�~Y�x�Gձ�+���a.��>�s���ooK$�w��V��l�:̬����׻�:�剅-�Tb�*�1cFL�����_Uͽ���jVؒߧ�>��cw�5�[|v��,����	� ��@�'q3<zx�� ����UIR5b��i�TE�˕�~EŬ���tt�m�,�g�*X��D[�_O�" D�؄��礌Xzޛ�q�9ٛ�U��A�-#zd�o�,&}�z�P0����ly��`����vL;ve�?�1�ؗC�;H��;K�ݯF+�v��L�;�~y�u�%���"������U��U�Ѱ@�ܸf��f&8:@��E#��8��Y��M&W�1~���˵��N��H�)��Lp�N}!Z�j`L ?j�ț��y\��|�!�[N�}xkiI���d�S��i[FɎ3�;���!Y��{�T�>2Y��d��SY�9oK���v45�]���o��OH�|��I���|g0)�<W+J��j����Bڝc�Sʺ�Ry'��d����Y*��=��wX�-�[��t^���*�UF���P�r���5�WԬ�fN�u��@TE�2y�G���W*~*���/��]���n���������]��	�����#���#sZ�bq�{7�E��ߵx�e-�2�8E��oc,ۜm�$��2���zL#�B�qTfŬA�Ĝ�|��)�u��+:�;&`�<%(P$�Nq��0H/�����ƺ7�;A1�3q�����W��>�-�`�[���܉`2[,�ۅg�Oκ"}Ă��߿��#x=5�ru�ޒ��@MM��V5���O5�8�_��0��ۊ���?��8ai�2����S�!���K��V0�)�n�Үz�O���Y��rK���󈇟����'��Ek:a����'���؆	��@�7��~�bBZ�@3ܡ���;�fL����dw��V�̍0@j�vh`�`��X� �>�.�ą�>� ߸�z(WV��D����)p�.���
-B��rO�v�F(��any=/�������4�j�b��'�=��OQ�X�#��F0܀*z��U�s��+�r�*L�߼� ���%����ի JI�WĊB����R����E����P�#�%�=J�S�W�5����t��m	�o����Sy��r�ץ*��0��"���ޱ����mOKO;��4z0�8x��5��X^�gZ˔J��̤���(��?����< �H����;��Gn��B���<�����g�P�� Q�΢P_�'9�b ��x	{�Tah^ �;ɘe�2��S�Gr6���z�Cc��+�W�w�y���ӛ��l(�lO�n#��Qۼh��(�z�$睠�D#̜F���e��7�'l��"��#r�^�VJ��FP�~��dh�����R�C��BD};.Qno��������FHY��jyl�իI���|��PtD�5{j 
M��@���Ie�)ċ�x���ŌWͰ �˽�CN��*[�
�3�ј&����i��!
Lb�(R�Z��Ӛ2�	U���*l����\���{6Is�G����L��d���؎�8#��64���D����Į�`!��E�����R³��5�	�C�P�ߏ�3�i7Ӱ3��`��H/ڠ�;���w���h� H���/B̈�1,i~�
�F��N*0W�=�AD��}\k�̎�DP�(��!�|F�Jn.�IA@���MV�ɼ[ۏ�H�d�������F0tm�=�g`\���+�=�M�=K��n؟K�><r%���o�2O���~j�f7A@@M���W�0ÖCQ,v(oГ�v�	m��el�8WgJ��v8{�t�k�1Ø��i�.+I-�E6�0ur��5�:T}~����	�����U�P�Z=]�]BJ&�1}7k3(�/��ui�:XSh%�;X"����.�h��I�����?q��ӝ&��N�=P��=��h�xeǌ�ʳvî>��P"	"����`������O�l(����\�v������?t1�a��)��(,"'פ��*��l�5��wE~;� ��s�w�#<�C�5��l/$�8�a��������m?Ę^��ق(�6�7�=bKM|�sѓ�6<�"�R�1�ߡ��9����Q�r�ԫo�i
��zW��}<��c��b�����G��Ё�a�n�^dq6y�4-�4�ue(�fzj�g �Kw���K��� �����E�����	Z�������S˨��l(1�
��X�$��yWA=���Ë|����c~�)�ƃ!V�����~���M댞"�,�����\;��:�_4���x9���+�c����k(�e�������p��F~��0�zՐ3""@�W�-����a�K�#�Ű�s��so�	�`�K�"����Ps͗�r��(�8`#!I�]w�Y����|�W^��m�$���&iԢ^�W>w2�YW��4����_�PZ��:R��-T��75�/S+��HB�$�W�	�ff�d���&�||B'E�;�>����7��G�y�۳����F��o�b��_�ԙ4��p�|���g�l��;-lo�K�|d'~�1j7���:u���;�7����Zf�s���q��]g�Zm���1Tܰ��x����%8�#:tP}Gk�0ʂ�*�0S�!ڧ��Y����=�ρG2��m,l�¬)�Co[��4��\�������Ut���&��W���RL�A�7M�E0��=ɶAd�W�&ɻ}�<������l�9<����u�"~6D��f��K]İWGU<��iV���{�	�p'����
�� B�R�j?�T<l�J�J�����y;f�m[���XQM���[ב����Ҙ|Q3qg�~�����}�G�� ~�&������{��m3��Wrm(i
z�:p9MV�E��<?�	A��..��ά�Ρ_��k�gR���	��	���	E�%ЃA�g8����HX �$7���8���D+d=��8�� y�w��� �U��ܻ��jV�C
�D�U܈��~?#�L�r-��-��ђZ}�''�d����L��(�Z��I{����4S���̐��u���ə�GڅS�U�,��׼�o������!+����H�e��B�g��(�U~2��;������>ئ=���:�����ۙ����(f�1�3:~c����Udp�;5���F߹�wc� .?���q��&&O쿱n
B_�Şq.�ո��D<�X�?"�n�B��&AS����!p�`״�p{��i����Ɩm�s ��o���j1+o�M��9n��,�嵠tV�Q�[�����u��\����|R���sN��Uyn[>L�Dj�����W�`3U�Y�A�����2�h�����E�c0O�����¸�,��Z�?)w��M=u�JY0JH@l���k�[R�>4Lkh��S%;����8���R��]�Q�/1�;W���k�󖁙5��x�����a�̮I���UM��c�:����y�T���ڟ�p�� �$!�}�,c/�z�Ռ&���-�Ȃl7*TI�|s�Cp�� �Ψ^o�j���@g��E�Ҭ�3�|�؉&�~���@�7���+��w@�Rd*���)78�-^�� N�K��,��d�|�zƔ-ڌ�]A)���'�]����{r;�R\��2QPiZ��?ք�f¬�ܔ�+� ��^}��U�B�ȫ��Y5ju��ŅK��3�1'R����!߽���K��G!��k)v5��vs\�3q���@�s�(�M^7GOt�y{e��f�3�̣+@I�M�Iũ�Y6��3����G*��!�GŨ|��b�#ZkO�D[+�Y��&�!����4S��=�ː��p�xC����m��Ec�i�};^������Q �I�� ����OP��C��O��d�&G�9@�u��{��C��4�1���-<��o����U������k��Ph�k���8o����Ҋ`vG�mCSg��������ۈ���j^�Z1�=i\2Z���޹(a��?�O(�G� C
[AVJbt���VB����؇�.e^xP'�5�OÆ�8����,�p��f8>���!63S��E�����@�)Ƴ��ۉ��d���׏&u�[9i�Fԯ�1������@�J�����+mgb�[��'��J�:(�vX�7��7��U�ʇ��-@I�� ,$�iVȁ��8�f��da���,�'*!k�����j{���*\`��p�W�>���*!�N�vhZ��=������cT��T��@e�Ek,���ىi� �i	��[$k�|�E�qi�sf���H�������g�x)�Μ�9�R����$�A�}��{�kaQ����[��U(S��G�A�����v5e�ד�n.6|h����Z��#ĮIlYQ�n�ʺ������
��|o��aov�$�S�8��&7"<3( �BX����08fh�5�P��^����C'4�&�<y1��KV���p
�#wF���JQ��*	�>A(�S5P�yw86�܈#Ϳ�v�Ѐc
����ôQF6�Z\.3L�:��x�ߘbP"w�FLr�����k����%�!��8x1� 6_r�d��(�@��1x'��Dj�: