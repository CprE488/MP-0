XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���b<���wC|,`|�jK@�:�G���	�$� ��4:d�V �pp`�<�]8������2/�$Z�k�X� G.0䵊~����~1_ �l�b��pP�F�����:�S�I���Gg&��fC�����	��c>���$ �i���+U�m4Q��?r�
�l���`��qu&�VͦO���hoiv|����$�����Zٖh�F�5p蓜È�m0	�Kr������j��ll�H�e�a�����}Εꑎ�,�ʲ`�gs@-�/��Q��(�p5�	®���n���;�O��L�s�:���_Ť�Oh^G��E͘�c�\YK��^T�x���^6�i;��&�;|0N��h�,+g1�Lm��f��IA�- 7w��!�k�qq�AV����煊Q��$�q��X�5�Ut�|��I�Vʮ⵻W"}-f���Xs�G��Ǳ���l�ϯ����h} _�_?��9D�p�����ǌ�$S��5BNn���;���h;$3��{g}` �r��� ٣A~+�?gנ�~z���r�@�0* ^��2d?UM�J�Xϳ���(SR�h��������-{��u�Y�06z������� ZN)	P�
Sh��#���p�����.��|��Δ&)��NR�����-i�ٌ8�W�k�oL���	�W�u����{�6���H�!|��\l�kM��bG���Dq��%�=�wq��L~VP9�I��sO2�U�����#>�����i���/\XlxVHYEB    6346    1790����e2�H��ݘ��!v�m�Ij�@�Up�����^�J�.��$�։H���!|�j�-��͡�G�J_��������Fl�B�_�1��9��<4�+cq�?E�$��Bh1}o����7�aI�g$�{�_�L��^��TyBa^�,sd@�n��1GkPRW����A�F�6^�@}4��~v�e�%��u��{M��z=��'֪<�tsx_�����$Ɖ%���`uB,�BG�����oH�Fi��fN;��i�D`_P�����i~}z�ϟ�'D�0{8��R���3�K�N�\'�1�K�u4�R6�Xl�O��n�%��a��)P��KXh]�ϸr�#"��],�1��6���=�������<�x�Ԑ��%d�c`���#��M9��X`{��GX,l~�/6��e��bA�O;�.YA=��q���Cl���v�y!б݋���gS;|0B�v�q�ár)a_4�ͤ+%v��{�,NyOyS�m��T��b� �[��k�u�`�vUR����p�sƈ�	���l�.�<�̮���F�P��_?i �3�e�P�/�������	�R���@9�$NOyp7>�[�J$��^WAc0��x����,�W��QJ��pI��Rj]�*��KÉ��	�d}������^�X���5��H1�R�b*�K�T��q��!E��q*}��NIJ��ݖi^GҢ�A�s ��{M��B�?�U�=f��.S�-% �
����)��[�C�u���琾ϴ&+Ѐ���e������'P���J���i�Y��#�Hx�~ֈKl�4��4{�~6?gEvI��n�C_%�{�y��]i���n��&�u6�v��a@�(��X���i}����0�h��)�<V߽ꚿ稟$��m���g<c�CƖ͡���	l�0���ӡ��/�߫|�\�5pc�@Z�4����Ϻ���G�"S��9S)��k-}���jgK�Wǒ&_1� �ew蕫��7��@��0��ev��A�����A�n��>���/�f����&�A���v K��:���'a�1�)���&M�uȈ���� ��u�	��IuE�+.�(�d;ז��ۑ
����~[~�#k�22)zi�Q�	��w�\�"�~��e6@����]s^;
&هC}�4Eqa�<H�t�5�J��;�D��
E�$�����s^�?I[F"��  2)�N2�<�����
�U���X4C���;ܗ�1�����;�q�Էޭ����%���(��{HH���n��_�H�zhFU�sz����,�HZ]��!-<�KA$�M���-t��.w��̅>� k=!�.�<j�G(^�P�ր�l��Xﲔ=���M�v��h�
�xy��۶ZG��G!��1D�����F�/�J��@�	�ʏ2s��G݌)��X�Saf5��\9�S:��=c �t��`��NM��|��9-&e΀a������<�eV|�k2�fb�{j�#}m:��{����kc��"��NLu�(��!��9l�-�£Y���M��ɧ������jI�R����S�/��Ԏ�L��C�E�Um�~SEGF��*���7&Ʈ��=I��r3T�)PhK����#E3&���6+�f���:���,�0�v*j��'�<��Zu�S�tr���^d�����[�2��g��|r��Aaz��	7jCRkX�5��'V�s�,�/9z��)w� �;�8��	jCRb2�[�O�H��)��XZ%懊�x\��nX�����-����wa=���d9k��� �	�M��a�U�X"��"s�oòmld�@�x�)qX��v�t�"���]4s	<���@�j;G�C��b�]a$˱��b�t��Q�2x�+�����qr̨��G��JE��Wo�� ���v긾��y�sAC�^��-��(��A�}�	���CRU4���/e��Zqy�ˮ\<N*�o������\��_)��m���Z�s觎��IL�.�~ZPs��m;}��:�WP7#>Gx�~��ݲKQ#������dJe��a%�F$�E��eGQ^X�A�	�S�K�ȑ��W�w���5ř�za�y�ɲ�f����\@�{�U2��Ǧh�~Ӝ�:�ly�d��5�o�*a��#���0V���a\����ؼ���}��3�ڵ�Q�mr�ɏҏ=��N����W�t2|�
�&>IR����v���g�.8i��}K��Z��f֔�rP�>]��B����<m�$8]^��8|6��bh:֢:6���*����~˲c��orP#�IC}!�c,��Ah�1؟�3K�&A���~�B4Z�Ϸ�?���͍���͠Qu�{Bȣx�\ld��S�	�*N�U��c7�7\ӕ������b��}��k���Y�"�(��s���>1�1���3�r�]�ѬŖ� ����	1��%����/؇��Լ\��$㸉��=B; �;������t1�W�I1�T��q֝���0�������@V�4�������-�����2Y#�u �-\i+��#�4�.��	D{���xRT�)���8x��cl�]N)�oS��r��F�
�:R��vE�������|�P��W�N~���q��WA��|��\Ї2,���D��e]#��>*p�
n��{�q�J���k����~c.f:h"���b ��^���]Z}��]8�Q-N)��o�#[rG�#v�@�S���W�^����ZRs�G���b��9�:7 [�ۆZ��� m�Z[DgY0�tr��h�RGp��5��>��+s�&nѕ�n�]��l�
��2%�%����M�#�:�\4V�Tm��"�g4�
"s�l�(����_*�h�BC�w?��#N�Dt�H!Ye�s%)��@F�	�>�Po*��ɲu_~F��Rs�欥Qx_}���&�xi|p�$�뗔}����?�/���%l��G�� $�1�b�
��!�D�\�Q �@������KB�ڥ� ��}�T]��o�i&��"�`�mo�B��e�Χ@��D��X��T��K��U����
_���x���N	��)��!��J<IJM
kA��@��|�C�ÝA�u�7i���")�3�c9ſD�P�j����op%��ߴE�=��� |E�9���� ����{s	�ԋ�H�$�Y�x����ڛ��e��kN�K�S�*Զ�����r�n/p�Ϊ/m���#��xZ�)CXG��`�q�����'B�c�Z߽oQ2�>�>*Gײ�/�b�p����J��ociw�G��DA�G5��|�g�7Z����02�9� ��1��,W\�j�k�S�q��#�O8��i�|/��9��N��R�������1��v�}u�]^K��;�>���_<� �[2԰���w��RZ�������=.�./�u٫����<^�M4~q��+��Q��/$�������e��=��n���������~i�D�`Y��&�O3m%-�2��)�9FPB6|l��FM���mw�9��#�b��Ot�2aiE�p	~��+S��*g��e��]�*շ��{�I&'���M��7�7�ɣ��vI�(�{��g��)��!�է[���^N�Zm��2]�Èʞ�0���6'��ޛ��r�(�~)e㬆?3��Ǚ�}���� ���M>B ��,%��`�o�eD~U���_�}3'��������5Ĕ�[�>!v�����_7��ږ��hW�z4z�*Tm��a���ަl��5�u�����O����<��2�XZ��֭_�"J57�kD6��8� Q6Vz�bրk"�(}l�%8��"7�@k�O��1�d�|W��V�B~�Oj��F�Me�ӵ=����HAe�l˯�)Ӏ�����Q�P?p<�Cz̫�
a�W!Hw)�h�9�0�V�k��q���~�n���(�wUc)�~g}.�"��W�5,��c�}�@qm�+���>��^��KcXi���d��s�5̑^�����&�ؤFB=Z,�~�xO/N�����	���*����	y��2�"�� �p���r	a��i#���	}t�͇F<� �m���R������K�i<G��҄��د e�u勽��r�����������D�hngpr!T��л��\�T���U	��&8��un��	Sb�y��t�Ey����u�p�aZ��F���"J|���z �����O�U�ٟ�E��Y��РK6
�^/��ԇA�@w+Z���(K1��X��u�>��Դ�\�>��.12�,&r�}+ϡuXq��!*���qߐ��4i)�8l�v$��V\76R70�=��jD*%4�lS�:E����5� ]n �Uo���k��K���ATЧk�` ^l����ɀ�8�"�8��j,I~�f9�C&����U��i\C��.;�5k�dg�� W���u�\(�r�o�ʖ(c�ޏoXܺy;�8W��^���
ԫ����kp@�\�v>�&׬���<|h��$������o	G����8	��
"�W��f��D7Ow��cd��񠂼������<��dJ�>Q��H�ӭު���v�nz��BSmha������A���/Q�7��8l�I���_���h:����X�Ecka����z��)H*�������s�ڒ"��7y�������-�a��*M�cD��ݩ@_��jG?���[JG��Mk��gQ�[���3�!�$-�����OoS�(�(c�Wi�D�6J�!��{:ģ;,�]ĺ�'���r����"��Cf��I K]*9�����y��J����B�[��́.*��.��2Qx�>y9����V~qz�����û�Of�4M�H/�.�x{1��u?��{��ɯ}��)���[N�)*}%텱7~+�*[]�U�7eiE�:�&�BeY)�+N�Z�;f����@�˟�Ka���DM.�"��}��V�*�<D��������`7�ve�(;>D	�`&�8������[r�r;�m���� ��m�<Krҍ�J���w��x����Q�Ǳ�X��ɤVFBL������EE����1�%R�HÁ!g�|���C��٨1A�[���C<Jx�v�yVpM��� ;�����e�v���M�A�I��l��L�u`�d(�����e�[)��h�]�Sh[���
{9)�����e�A����pF�E��"(ȄE7��Vp=*�� ��[8i�󴡞K���e2��}yJX���`\S`�hJ#��B+�|W+&`;�fpm[#�(L����h�#�6�~zY�^Z�Sg�y�����8h���� +1�d��k͓�gP�A��)�;(8e�ЭA	�����	�d���V�S)���䘕Ȗ"ԣ�R����U��W�q�k�@kE0;�U���O)���T�R���=l��<�rwX�&��J����J�@H���e��V�6�sr�[��J��;0�7�r���9)o4B����Xŏ$?�%�c���Ly(��v���o��A�o{F2���M^���nz���ڃ�^����� PD'o=��~}L�w���#���4���ƖP��B0Z�>Yv��z�e#��#N��DƷS���;���J�B��+@ob�(�@�6��t��Q�@��(��C<�E�[�iSM�?X���}��x� ���b�ء#49�|�s�KǕN���O�@��[ljj�y�3(��e�b�ibw�2�3$�h�`�r�S����A��C~b+1�v8X�L"���	�"\ %3�`>3�7|Ƈ��F�%z}����Nl�/ҁ��h[��4D��p�p�"��D���G�$�Ud�"2S�އSR�RɉՙzىHv�9P�V8d���^n^�tq�3�~��
ʖ@oF��@|9�!�X�Շt'Q