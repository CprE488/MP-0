XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��n���$]_�����WO-�,� �۹te�z>�Ȉ�������"��L�A���g@|�up�O5	Gl%~�JJ�9Ǹ�^����8o@0d�5����E�V����O7ow�U�|�2aCS�~�R��$�$k��0�,����8��t6iY�m8����)�XGI-5� +Ζ_�d�۠����R�,��vT��<X��⻣�i^=����t��>BW�(�_:���2��Dc�bEc6�-K\L)h��.\���6�[������v�r��|���Q�
|�F�PXL��n�D^�yw�չ�U��)0���e:;���u�̀J�p sV���̤$<o?�cN!C��zO�A��<yЧ<H�?2�n�q�ypԀ`�4>��<г�!�	-o��K���z�}��t�����]�ѕQ<�@E�g�/���0a0�&���R���ma�`5�eg��ZѾQ���G�S��eÁ�G���8�PtT��Yrw�R������HZ^z�O���RB.9Kh�t����C,�O�8 |=3Q"2ǩHG�^D2{��w}ӽG��$"|��WI��XՄ��A*��+r������!GO�_Ç��![[c$�>���O��V<��i$�}b�k/�5�K;O���ȶq�.ĸ��_k|s_�`�����V�Ů�C��#Bc�Y�/�+U7j(R/uE��#b�o~��N��j�J�o>��e����j$�A�_��<M�� ��e��,��Y�.�w��D�����j�w�q�XlxVHYEB    42ae    1110��_&7���@���ʊ0����M^Mb�w'_�	�pXy�|-�aM*\)�PxA��ˉf�M����n�l0}A�}����9�$r�˝�ʹ��D� 	@:���K��]�����HO���1�q
wlq|��Qr`��YC�NJ�Q�$���a�W�^1��#�<3�pP��A�j�-�}WB����RX\�9��7�F�j��_�u���e��+�R��Դ;��.�� 8C���-o�$�|����٠�{uL!�{����r�Sdy�-�K~3)�5Cw�l �b���rO����r���ULe��9h�·�x7:���Q�/��h�\�7]���i���tl(����}��P�+�y
�O܉����!,_�j�c��?Ɏ�32��,�
E�55)W~d%۩^,1������kH���>/1� ��x�?꽍�����?�ǃ��\[|n�ba$�������'Oc�t�j�;��ڥ}Y-�@U��IP�ĕ���
��^�E���_�J_jzl��WKd��:��b�����0��}켅��܎<�D�����m��}J��և1�]�͎�ڜ}K��G,68-9��K<s��R����zd��u,-|W��]*�x�2;��Hɾ���U��?�1G����f^� ���|b��䰯���+�%�����<��Q$�F���*J e��DU�y-�Ϸ���w�߆���h���-�q�i��߁-�f^�B���YƢ��I�\E�ue�t�Z�.�A�ͼN�=����91W��X8$��9��b�"ܓ���+!yn��F�����	iFQ��£��'�b�8��'ʋ�F��pX�ԙI�f�չ�@F1���6�)S�\�)�\����-�~A�M��6����@٬j=~u[ݨwh5v�Q2�u�-K��@�<��k���"��%9�^"���HX�.�1U��ۉ��k��g�X]%`����>�����^U��G�[��c`<�>^huMI�F���r`�w�fpbi1s�����x���}���^!u<h�~��#zL 6�"l'�V'�Z2��n �>�IB��:��N�/�)���.X�+m$�^P��yMZ ��m����`qr�k%���|,SE� ����-�tC�, �4����~j�����C����v�ˤ|��)����ceU����pmЪ#�r����E�<:Tk�~pn�/��,�����i��#^F���u%��&H�������F<��v��1�/�C �4���Ub�*2�8���E�7����C08)��	�"�Z�5�����T�A����$Mٺ����kʝ6q�����4�B�u
4�Z��c�6�9r�a��-M�N�����c%��`�
7� �H�~�i�\=(�q)����I�ya,������S�ߒ���>fN��k�0�ז�?�"�o����hJ���
6l:��k��b����bZ�e�hQ!Cn����[��왝�n�>h83ߍ���W��>z�<I4��x��1x����pݿ��
asS\R�>��2l^\7���� A�7�o�"���%��|�q>��7JN�
�v�e��`�f�_g��;� ��%����B�Z���w�ŷ �g&#uNbE��l�L��vt�Bόʈ�]��-�x+&xni�a4���y\ɲJ�K�Jy�Ճ�E�������jX�"9M���>V?��Y��~�vV{H֭X�����Eyۋ�GSB;��;�.�l�m��l\e�~m�Q��֛��
,�tF~`����V��B�9�p�.W��=�mk;T����ڲ? 9DV�H� �o��%c������#V7fg8�J���4� р�w[+�bU��:f2��2 7��)������P�i���n�"rc���֬yWt�O���,ί�=�~S#~a�*��G!�O=������:�͎�ކH�5�� Mp��v��Ֆ�U�������&ǅ:�P�q���*gk6*��$���ΒJ:
^z�����/��Ƹ3�h�!W߰�"�||5����G�=��M"9Xx�`B�r�c7���*�zmb�����׀��G>ABl4+�ލ�I�a:��0'�/Ҳ�fo4<1I�M!��.@)�&�V 7�� .����g'�1��q�Hs���!�Z:�A97�eYM�w4��|���)+m�g��l"�N+�ʕ���:@��
/H�n�L�>'��Yr)	kg/���0��O<4P�sY�h!L秂Q 1��a`���Er�e�C|����]�y�nޫ�)r��QH�9�^�Q�L��b�)���(#�~9q��͋ū!6���#R�������E�I���f7��ři�(O#�'4h<w�l���8�X �뜨���k#�����6�Y�L�<4�&\�<<��[/6��f};Oց���UA���j�q�?O�L/9�}�6��u5@s���7��%E�����R� <�#���Ů�x�գU��Ie�s�C�u�^��}	��a����9�3]p���52�q5�,������^�y�n�s�fO�T���?�
���ڤo-\�e���w�C����^BM_ʕ`�l�m�2NY�p�gX����=����{u1�j��hI��FP� y*.��h������+ͨ���ڹ��m�S���M�E��<jW��-�o�����u,�k�N�3-ߨ73�b����zu��<R��5X$3Z��)^�1��.xc�Wc�G�J��q�\�XO&�	:sM����%|l-�� �.�*5�5���匫�p���k�G�Q��:�kӗ�O�Yv⁪����X�{No��5����vY��l��K�`Q��	�"������n�Q�L/<1���С`�s# ���`�	Շ�+�F�<������Iow��^ĄtC��4"��P���r+<Q�i����:�|�X]�ĈAk7\�z�|).e_?3�N�����?7�@)>��곰}Ve�_�+��p?�t��I��s�5��9�oQM{o��w�q�T{̕�:s�J�*k�`��DmH�����\��|jtbp�������Z����Pn��+[i�ԕO�R�0\�\��J:F����[S2� ���G���&��*~$��l2�wlI���>�qT�o�z��$������̫Au��f�)(h�Q���S�>��-�m�4��E϶���6�~����^�0�jY'�4u_��§m�7���q�L?����Y����8�2Ors������龟9�����&f�ub��x2FG94���_
�@fg;���<~t��[?�c$s�sɷ4t��#��n'_\Gد6p��IX�2؉�Ɔʞ�4���N�V�d��
��1z�3�Z���Ҽ[ZSI�'</�<:� ��`&�����I�[7��HO#�!`/���V>��`�YP�{,��s�
\�<3)y�%�;"���5a7�p��C�CZ��٥�tp�+�Xcʙ�Gm���[9w�$P�M���a��<�V7�M�-�J��z��v���������QJ`k_�8�%ւ(Ȫ䋅��~�C`r�߫���/��kALɕ�Vb��T�Q
��$��F��ӃC��`�q�5���)\Y6�����D���J`��Z�9��xl��y�o�rT�쇮�G��o�noj����w��h���a|i+���>����Lu��Q �)�D�7	�,�p���O��\.g��3���ڜ�_�BJ�6�G(��㧩��܂�����M"��H��-�X5��τNMT�s�qPX_�w�����	�u��-䟹���(g;~N�	�Y#H��z�DO��� �}^w��C��{UE����
ֆ�|��c�W�`r�"�����hp2�و�,��n���R n_�9<���?���z�$��-�So�����^��o�[��3LJ"��Wi����o�/g���7��c7����1�	��Pk!�,�ǫ=�*��R�v�h�hv�(S��"*9���1�Ji�⩛'G:���4Ѯj��&j4��#v
D���u�wt�3c�&0������E'���I�d13�T;��L
	:��kǭV�P	�y*�خ{�_,�Y�)�9���.��LX��5�#�4��&�/���7ј&9!�81w�r��-��;*���WM6(��".
,�
`~��	U���]��r��5 PLE61��@D�	�+(&��%>���_�B�����|��?7�1ޠ���*�e"kG��xDP��p��]�;9W?RU�G~�V�