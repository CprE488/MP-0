XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[1�Z"$����i���Zhh%�t�����|����D��:d����|�t�9�0ם�����-�i~e������V��E�9�q��Jd��td-���JyQ�m�MT��P� ���뎗b�m�~2x�n~���q��]GK��~�I�m�)�0���C���X��oi�xo8��E�����yǔcӡ(6oJޠΜ��RmX�� ���7�%���*��PY��ht��P����M�.U1�[�w0G�r��s��4���>A���f塸��!���@.�졿	�ד7�+��e��K�����9̈��¶j�v��F��$>[���9�������"1����]�!Vblh r��p.�v���n	�����,���8�^�J6��T�t7`$��[ywo2�aK���f�M��V`���L��#@�U��/��z�*�L:���[��wX������A��:f1Qim�H�N�c �_�!�R^�Q+��a�cG|`x�`*9���)*���}-��m�c�C~��XF�ި� ��4�$���!`�W*�_]���X��%;^Z�yM~*��A/K�ڠQ���i���Ui���+@s� �]"�4��~ l�Zei�AGXWXDcaS���͹-��P�ި)�K]!�����.WA��rp�*�ԍ�Sp��F@��(^j�8�s�9|���.�>gH'pǷ�C/8ŁS:��TI�N�U�3^-��7�@�NgЎ�{���KD�,L���UA����XlxVHYEB     f6d     6f0��~�0XE{���|}P%0m>z9J�ܰk�J@�m���ͬ�F�L��gpm��v\�P��2Mf����R��.��oъ�a8�<R���%1�z֭��Ar�c��&�j�m���]�\�aKH���3 5T{��J��#�.)��F�hO����@��%�bTF~W1j�E$%l4�_���>�&É���n�����"*�[�S_�MqÇ��J�4���o
C�Q�W����^pF�Ӭ�u�ݺ��6���XH*w
!i�S����o&�*"��r�Ol��ꖹ���p׫��8�z����ڤn�H-��e�r�f�r����b��f��j����:@��������Ƶt��0��m�	T��2E�<o��2PqLv@@/���2�p�1�܀�mGԂ��~Xs64�< {�Пp����~��E/�@�h�9l���g�33h�3ki�e�o�$6����ʗez��h*�s֘1EC��#�~sX_� rD=�ぜD&j*�k`�����H��V	ի�pYИ�})ґ�̿�"���1âO18�^e����6*�GHE��N�1�M7~�4v9	Bb֭.�<2iW�͟+>w߾�(@����	:�����Rc�w�"d������i�⫞B笍�x�n�4	��bs(Lp)eW�Քrw�j�Z�����^�f�Ur�#��a	�k$me�)�3t�P9g �5)��;G�#���xQ�9�T([5�dߎ"�qi�wߴ�E�T�B�r�(o�]�r�ߵ�,1Y�`�02 ��v7�[S�I\��떬4e��e��Ef �H�c�:�g�V�UMaC3$*�D�h��FZH*�,���c4:�A����T�p�=pc�d�8Vh%���'�SM�� ��T� F�����"XNQ���!{�%c[q�d✛�VY�2�CL��y%Z���s��X����B��ʒ�=��D��}���0����U��������H��d���>m �h��C���-�ѓm�H�6�~�U�:_QQ�w�jؙ�%�twc�����7�S~�%�A`4	 �sb�,EK�U��I��:�	)/mt�l@�a��ny))�O�Z�q�"���*�bO��M��<ԏ����d�b�FX�B�;z ��̷�3N��16ˣ�VB]`�NZ΋��>hcϰ��,7k7�`O�%�̃�����'C(��&�<�x�duy"�2�$ī�ŕ��b����U�����qUU����ױ���R����W�՝ .�O�C�1�^
������ĳ@�㩈O�=ɩ�'(sV��E��.�3껇��I�;���Q�)��O2�5X�ѫP�z��焐��'Rn"Ι)b= �z9�ۏ�m�"�E�xA�O������L���K�����=�T���>��cX�I�"3,� ��<A����IsYAp�!K�C���7\�)�B��2f�z�� ����A)��'�t���$I=�G�`��Y��@��?tw�!��5 �*����f�z��G$'�r{��H����8~F!\��My��3L���c���{p��aQ���		��=�0��+��8W�
�Y��6@�K�噏��8;�`�{֘;�bx�{�u�AG�m�. ����'�=Ъ���?��
�����x=������n�}c;ya��9��ێ�څ�U=�S�N��\�Z�]�ڄ�#�g�&:T���q�䣶�c����x�|��Td-�4�)��3��8�I��:v�D����T���cz�K����